`timescale 1ns/1ns

`include "common_types.vh"
import common_types_pkg::*;
`include "multiplier_if.vh"

// Wallace Tree Multiplier
// Pipelined, every 2 stages

module multiplier (
    input logic clk, nrst,
    multiplier_if.mult multiplier_if
);

logic weight_0_0;
logic [1:0] weight_0_1;
logic [2:0] weight_0_2;
logic [3:0] weight_0_3;
logic [4:0] weight_0_4;
logic [5:0] weight_0_5;
logic [6:0] weight_0_6;
logic [7:0] weight_0_7;
logic [8:0] weight_0_8;
logic [9:0] weight_0_9;
logic [10:0] weight_0_10;
logic [11:0] weight_0_11;
logic [12:0] weight_0_12;
logic [13:0] weight_0_13;
logic [14:0] weight_0_14;
logic [15:0] weight_0_15;
logic [16:0] weight_0_16;
logic [17:0] weight_0_17;
logic [18:0] weight_0_18;
logic [19:0] weight_0_19;
logic [20:0] weight_0_20;
logic [21:0] weight_0_21;
logic [22:0] weight_0_22;
logic [23:0] weight_0_23;
logic [24:0] weight_0_24;
logic [25:0] weight_0_25;
logic [26:0] weight_0_26;
logic [27:0] weight_0_27;
logic [28:0] weight_0_28;
logic [29:0] weight_0_29;
logic [30:0] weight_0_30;
logic [31:0] weight_0_31;
logic [30:0] weight_0_32;
logic [29:0] weight_0_33;
logic [28:0] weight_0_34;
logic [27:0] weight_0_35;
logic [26:0] weight_0_36;
logic [25:0] weight_0_37;
logic [24:0] weight_0_38;
logic [23:0] weight_0_39;
logic [22:0] weight_0_40;
logic [21:0] weight_0_41;
logic [20:0] weight_0_42;
logic [19:0] weight_0_43;
logic [18:0] weight_0_44;
logic [17:0] weight_0_45;
logic [16:0] weight_0_46;
logic [15:0] weight_0_47;
logic [14:0] weight_0_48;
logic [13:0] weight_0_49;
logic [12:0] weight_0_50;
logic [11:0] weight_0_51;
logic [10:0] weight_0_52;
logic [9:0] weight_0_53;
logic [8:0] weight_0_54;
logic [7:0] weight_0_55;
logic [6:0] weight_0_56;
logic [5:0] weight_0_57;
logic [4:0] weight_0_58;
logic [3:0] weight_0_59;
logic [2:0] weight_0_60;
logic [1:0] weight_0_61;
logic weight_0_62;
logic [31:0] a, b;

always_comb begin
    a = multiplier_if.a;
    b = multiplier_if.b;

    // If negative, convert to positive
    if (multiplier_if.is_signed_a) begin
        a = multiplier_if.a[31] ? (~multiplier_if.a + 1) : multiplier_if.a;
    end
    if (multiplier_if.is_signed_b) begin
        b = multiplier_if.b[31] ? (~multiplier_if.b + 1) : multiplier_if.b;
    end
end

assign weight_0_0 = a[0] & b[0];
assign weight_0_1[0] = a[0] & b[1];
assign weight_0_1[1] = a[1] & b[0];
assign weight_0_2[0] = a[0] & b[2];
assign weight_0_2[1] = a[1] & b[1];
assign weight_0_2[2] = a[2] & b[0];
assign weight_0_3[0] = a[0] & b[3];
assign weight_0_3[1] = a[1] & b[2];
assign weight_0_3[2] = a[2] & b[1];
assign weight_0_3[3] = a[3] & b[0];
assign weight_0_4[0] = a[0] & b[4];
assign weight_0_4[1] = a[1] & b[3];
assign weight_0_4[2] = a[2] & b[2];
assign weight_0_4[3] = a[3] & b[1];
assign weight_0_4[4] = a[4] & b[0];
assign weight_0_5[0] = a[0] & b[5];
assign weight_0_5[1] = a[1] & b[4];
assign weight_0_5[2] = a[2] & b[3];
assign weight_0_5[3] = a[3] & b[2];
assign weight_0_5[4] = a[4] & b[1];
assign weight_0_5[5] = a[5] & b[0];
assign weight_0_6[0] = a[0] & b[6];
assign weight_0_6[1] = a[1] & b[5];
assign weight_0_6[2] = a[2] & b[4];
assign weight_0_6[3] = a[3] & b[3];
assign weight_0_6[4] = a[4] & b[2];
assign weight_0_6[5] = a[5] & b[1];
assign weight_0_6[6] = a[6] & b[0];
assign weight_0_7[0] = a[0] & b[7];
assign weight_0_7[1] = a[1] & b[6];
assign weight_0_7[2] = a[2] & b[5];
assign weight_0_7[3] = a[3] & b[4];
assign weight_0_7[4] = a[4] & b[3];
assign weight_0_7[5] = a[5] & b[2];
assign weight_0_7[6] = a[6] & b[1];
assign weight_0_7[7] = a[7] & b[0];
assign weight_0_8[0] = a[0] & b[8];
assign weight_0_8[1] = a[1] & b[7];
assign weight_0_8[2] = a[2] & b[6];
assign weight_0_8[3] = a[3] & b[5];
assign weight_0_8[4] = a[4] & b[4];
assign weight_0_8[5] = a[5] & b[3];
assign weight_0_8[6] = a[6] & b[2];
assign weight_0_8[7] = a[7] & b[1];
assign weight_0_8[8] = a[8] & b[0];
assign weight_0_9[0] = a[0] & b[9];
assign weight_0_9[1] = a[1] & b[8];
assign weight_0_9[2] = a[2] & b[7];
assign weight_0_9[3] = a[3] & b[6];
assign weight_0_9[4] = a[4] & b[5];
assign weight_0_9[5] = a[5] & b[4];
assign weight_0_9[6] = a[6] & b[3];
assign weight_0_9[7] = a[7] & b[2];
assign weight_0_9[8] = a[8] & b[1];
assign weight_0_9[9] = a[9] & b[0];
assign weight_0_10[0] = a[0] & b[10];
assign weight_0_10[1] = a[1] & b[9];
assign weight_0_10[2] = a[2] & b[8];
assign weight_0_10[3] = a[3] & b[7];
assign weight_0_10[4] = a[4] & b[6];
assign weight_0_10[5] = a[5] & b[5];
assign weight_0_10[6] = a[6] & b[4];
assign weight_0_10[7] = a[7] & b[3];
assign weight_0_10[8] = a[8] & b[2];
assign weight_0_10[9] = a[9] & b[1];
assign weight_0_10[10] = a[10] & b[0];
assign weight_0_11[0] = a[0] & b[11];
assign weight_0_11[1] = a[1] & b[10];
assign weight_0_11[2] = a[2] & b[9];
assign weight_0_11[3] = a[3] & b[8];
assign weight_0_11[4] = a[4] & b[7];
assign weight_0_11[5] = a[5] & b[6];
assign weight_0_11[6] = a[6] & b[5];
assign weight_0_11[7] = a[7] & b[4];
assign weight_0_11[8] = a[8] & b[3];
assign weight_0_11[9] = a[9] & b[2];
assign weight_0_11[10] = a[10] & b[1];
assign weight_0_11[11] = a[11] & b[0];
assign weight_0_12[0] = a[0] & b[12];
assign weight_0_12[1] = a[1] & b[11];
assign weight_0_12[2] = a[2] & b[10];
assign weight_0_12[3] = a[3] & b[9];
assign weight_0_12[4] = a[4] & b[8];
assign weight_0_12[5] = a[5] & b[7];
assign weight_0_12[6] = a[6] & b[6];
assign weight_0_12[7] = a[7] & b[5];
assign weight_0_12[8] = a[8] & b[4];
assign weight_0_12[9] = a[9] & b[3];
assign weight_0_12[10] = a[10] & b[2];
assign weight_0_12[11] = a[11] & b[1];
assign weight_0_12[12] = a[12] & b[0];
assign weight_0_13[0] = a[0] & b[13];
assign weight_0_13[1] = a[1] & b[12];
assign weight_0_13[2] = a[2] & b[11];
assign weight_0_13[3] = a[3] & b[10];
assign weight_0_13[4] = a[4] & b[9];
assign weight_0_13[5] = a[5] & b[8];
assign weight_0_13[6] = a[6] & b[7];
assign weight_0_13[7] = a[7] & b[6];
assign weight_0_13[8] = a[8] & b[5];
assign weight_0_13[9] = a[9] & b[4];
assign weight_0_13[10] = a[10] & b[3];
assign weight_0_13[11] = a[11] & b[2];
assign weight_0_13[12] = a[12] & b[1];
assign weight_0_13[13] = a[13] & b[0];
assign weight_0_14[0] = a[0] & b[14];
assign weight_0_14[1] = a[1] & b[13];
assign weight_0_14[2] = a[2] & b[12];
assign weight_0_14[3] = a[3] & b[11];
assign weight_0_14[4] = a[4] & b[10];
assign weight_0_14[5] = a[5] & b[9];
assign weight_0_14[6] = a[6] & b[8];
assign weight_0_14[7] = a[7] & b[7];
assign weight_0_14[8] = a[8] & b[6];
assign weight_0_14[9] = a[9] & b[5];
assign weight_0_14[10] = a[10] & b[4];
assign weight_0_14[11] = a[11] & b[3];
assign weight_0_14[12] = a[12] & b[2];
assign weight_0_14[13] = a[13] & b[1];
assign weight_0_14[14] = a[14] & b[0];
assign weight_0_15[0] = a[0] & b[15];
assign weight_0_15[1] = a[1] & b[14];
assign weight_0_15[2] = a[2] & b[13];
assign weight_0_15[3] = a[3] & b[12];
assign weight_0_15[4] = a[4] & b[11];
assign weight_0_15[5] = a[5] & b[10];
assign weight_0_15[6] = a[6] & b[9];
assign weight_0_15[7] = a[7] & b[8];
assign weight_0_15[8] = a[8] & b[7];
assign weight_0_15[9] = a[9] & b[6];
assign weight_0_15[10] = a[10] & b[5];
assign weight_0_15[11] = a[11] & b[4];
assign weight_0_15[12] = a[12] & b[3];
assign weight_0_15[13] = a[13] & b[2];
assign weight_0_15[14] = a[14] & b[1];
assign weight_0_15[15] = a[15] & b[0];
assign weight_0_16[0] = a[0] & b[16];
assign weight_0_16[1] = a[1] & b[15];
assign weight_0_16[2] = a[2] & b[14];
assign weight_0_16[3] = a[3] & b[13];
assign weight_0_16[4] = a[4] & b[12];
assign weight_0_16[5] = a[5] & b[11];
assign weight_0_16[6] = a[6] & b[10];
assign weight_0_16[7] = a[7] & b[9];
assign weight_0_16[8] = a[8] & b[8];
assign weight_0_16[9] = a[9] & b[7];
assign weight_0_16[10] = a[10] & b[6];
assign weight_0_16[11] = a[11] & b[5];
assign weight_0_16[12] = a[12] & b[4];
assign weight_0_16[13] = a[13] & b[3];
assign weight_0_16[14] = a[14] & b[2];
assign weight_0_16[15] = a[15] & b[1];
assign weight_0_16[16] = a[16] & b[0];
assign weight_0_17[0] = a[0] & b[17];
assign weight_0_17[1] = a[1] & b[16];
assign weight_0_17[2] = a[2] & b[15];
assign weight_0_17[3] = a[3] & b[14];
assign weight_0_17[4] = a[4] & b[13];
assign weight_0_17[5] = a[5] & b[12];
assign weight_0_17[6] = a[6] & b[11];
assign weight_0_17[7] = a[7] & b[10];
assign weight_0_17[8] = a[8] & b[9];
assign weight_0_17[9] = a[9] & b[8];
assign weight_0_17[10] = a[10] & b[7];
assign weight_0_17[11] = a[11] & b[6];
assign weight_0_17[12] = a[12] & b[5];
assign weight_0_17[13] = a[13] & b[4];
assign weight_0_17[14] = a[14] & b[3];
assign weight_0_17[15] = a[15] & b[2];
assign weight_0_17[16] = a[16] & b[1];
assign weight_0_17[17] = a[17] & b[0];
assign weight_0_18[0] = a[0] & b[18];
assign weight_0_18[1] = a[1] & b[17];
assign weight_0_18[2] = a[2] & b[16];
assign weight_0_18[3] = a[3] & b[15];
assign weight_0_18[4] = a[4] & b[14];
assign weight_0_18[5] = a[5] & b[13];
assign weight_0_18[6] = a[6] & b[12];
assign weight_0_18[7] = a[7] & b[11];
assign weight_0_18[8] = a[8] & b[10];
assign weight_0_18[9] = a[9] & b[9];
assign weight_0_18[10] = a[10] & b[8];
assign weight_0_18[11] = a[11] & b[7];
assign weight_0_18[12] = a[12] & b[6];
assign weight_0_18[13] = a[13] & b[5];
assign weight_0_18[14] = a[14] & b[4];
assign weight_0_18[15] = a[15] & b[3];
assign weight_0_18[16] = a[16] & b[2];
assign weight_0_18[17] = a[17] & b[1];
assign weight_0_18[18] = a[18] & b[0];
assign weight_0_19[0] = a[0] & b[19];
assign weight_0_19[1] = a[1] & b[18];
assign weight_0_19[2] = a[2] & b[17];
assign weight_0_19[3] = a[3] & b[16];
assign weight_0_19[4] = a[4] & b[15];
assign weight_0_19[5] = a[5] & b[14];
assign weight_0_19[6] = a[6] & b[13];
assign weight_0_19[7] = a[7] & b[12];
assign weight_0_19[8] = a[8] & b[11];
assign weight_0_19[9] = a[9] & b[10];
assign weight_0_19[10] = a[10] & b[9];
assign weight_0_19[11] = a[11] & b[8];
assign weight_0_19[12] = a[12] & b[7];
assign weight_0_19[13] = a[13] & b[6];
assign weight_0_19[14] = a[14] & b[5];
assign weight_0_19[15] = a[15] & b[4];
assign weight_0_19[16] = a[16] & b[3];
assign weight_0_19[17] = a[17] & b[2];
assign weight_0_19[18] = a[18] & b[1];
assign weight_0_19[19] = a[19] & b[0];
assign weight_0_20[0] = a[0] & b[20];
assign weight_0_20[1] = a[1] & b[19];
assign weight_0_20[2] = a[2] & b[18];
assign weight_0_20[3] = a[3] & b[17];
assign weight_0_20[4] = a[4] & b[16];
assign weight_0_20[5] = a[5] & b[15];
assign weight_0_20[6] = a[6] & b[14];
assign weight_0_20[7] = a[7] & b[13];
assign weight_0_20[8] = a[8] & b[12];
assign weight_0_20[9] = a[9] & b[11];
assign weight_0_20[10] = a[10] & b[10];
assign weight_0_20[11] = a[11] & b[9];
assign weight_0_20[12] = a[12] & b[8];
assign weight_0_20[13] = a[13] & b[7];
assign weight_0_20[14] = a[14] & b[6];
assign weight_0_20[15] = a[15] & b[5];
assign weight_0_20[16] = a[16] & b[4];
assign weight_0_20[17] = a[17] & b[3];
assign weight_0_20[18] = a[18] & b[2];
assign weight_0_20[19] = a[19] & b[1];
assign weight_0_20[20] = a[20] & b[0];
assign weight_0_21[0] = a[0] & b[21];
assign weight_0_21[1] = a[1] & b[20];
assign weight_0_21[2] = a[2] & b[19];
assign weight_0_21[3] = a[3] & b[18];
assign weight_0_21[4] = a[4] & b[17];
assign weight_0_21[5] = a[5] & b[16];
assign weight_0_21[6] = a[6] & b[15];
assign weight_0_21[7] = a[7] & b[14];
assign weight_0_21[8] = a[8] & b[13];
assign weight_0_21[9] = a[9] & b[12];
assign weight_0_21[10] = a[10] & b[11];
assign weight_0_21[11] = a[11] & b[10];
assign weight_0_21[12] = a[12] & b[9];
assign weight_0_21[13] = a[13] & b[8];
assign weight_0_21[14] = a[14] & b[7];
assign weight_0_21[15] = a[15] & b[6];
assign weight_0_21[16] = a[16] & b[5];
assign weight_0_21[17] = a[17] & b[4];
assign weight_0_21[18] = a[18] & b[3];
assign weight_0_21[19] = a[19] & b[2];
assign weight_0_21[20] = a[20] & b[1];
assign weight_0_21[21] = a[21] & b[0];
assign weight_0_22[0] = a[0] & b[22];
assign weight_0_22[1] = a[1] & b[21];
assign weight_0_22[2] = a[2] & b[20];
assign weight_0_22[3] = a[3] & b[19];
assign weight_0_22[4] = a[4] & b[18];
assign weight_0_22[5] = a[5] & b[17];
assign weight_0_22[6] = a[6] & b[16];
assign weight_0_22[7] = a[7] & b[15];
assign weight_0_22[8] = a[8] & b[14];
assign weight_0_22[9] = a[9] & b[13];
assign weight_0_22[10] = a[10] & b[12];
assign weight_0_22[11] = a[11] & b[11];
assign weight_0_22[12] = a[12] & b[10];
assign weight_0_22[13] = a[13] & b[9];
assign weight_0_22[14] = a[14] & b[8];
assign weight_0_22[15] = a[15] & b[7];
assign weight_0_22[16] = a[16] & b[6];
assign weight_0_22[17] = a[17] & b[5];
assign weight_0_22[18] = a[18] & b[4];
assign weight_0_22[19] = a[19] & b[3];
assign weight_0_22[20] = a[20] & b[2];
assign weight_0_22[21] = a[21] & b[1];
assign weight_0_22[22] = a[22] & b[0];
assign weight_0_23[0] = a[0] & b[23];
assign weight_0_23[1] = a[1] & b[22];
assign weight_0_23[2] = a[2] & b[21];
assign weight_0_23[3] = a[3] & b[20];
assign weight_0_23[4] = a[4] & b[19];
assign weight_0_23[5] = a[5] & b[18];
assign weight_0_23[6] = a[6] & b[17];
assign weight_0_23[7] = a[7] & b[16];
assign weight_0_23[8] = a[8] & b[15];
assign weight_0_23[9] = a[9] & b[14];
assign weight_0_23[10] = a[10] & b[13];
assign weight_0_23[11] = a[11] & b[12];
assign weight_0_23[12] = a[12] & b[11];
assign weight_0_23[13] = a[13] & b[10];
assign weight_0_23[14] = a[14] & b[9];
assign weight_0_23[15] = a[15] & b[8];
assign weight_0_23[16] = a[16] & b[7];
assign weight_0_23[17] = a[17] & b[6];
assign weight_0_23[18] = a[18] & b[5];
assign weight_0_23[19] = a[19] & b[4];
assign weight_0_23[20] = a[20] & b[3];
assign weight_0_23[21] = a[21] & b[2];
assign weight_0_23[22] = a[22] & b[1];
assign weight_0_23[23] = a[23] & b[0];
assign weight_0_24[0] = a[0] & b[24];
assign weight_0_24[1] = a[1] & b[23];
assign weight_0_24[2] = a[2] & b[22];
assign weight_0_24[3] = a[3] & b[21];
assign weight_0_24[4] = a[4] & b[20];
assign weight_0_24[5] = a[5] & b[19];
assign weight_0_24[6] = a[6] & b[18];
assign weight_0_24[7] = a[7] & b[17];
assign weight_0_24[8] = a[8] & b[16];
assign weight_0_24[9] = a[9] & b[15];
assign weight_0_24[10] = a[10] & b[14];
assign weight_0_24[11] = a[11] & b[13];
assign weight_0_24[12] = a[12] & b[12];
assign weight_0_24[13] = a[13] & b[11];
assign weight_0_24[14] = a[14] & b[10];
assign weight_0_24[15] = a[15] & b[9];
assign weight_0_24[16] = a[16] & b[8];
assign weight_0_24[17] = a[17] & b[7];
assign weight_0_24[18] = a[18] & b[6];
assign weight_0_24[19] = a[19] & b[5];
assign weight_0_24[20] = a[20] & b[4];
assign weight_0_24[21] = a[21] & b[3];
assign weight_0_24[22] = a[22] & b[2];
assign weight_0_24[23] = a[23] & b[1];
assign weight_0_24[24] = a[24] & b[0];
assign weight_0_25[0] = a[0] & b[25];
assign weight_0_25[1] = a[1] & b[24];
assign weight_0_25[2] = a[2] & b[23];
assign weight_0_25[3] = a[3] & b[22];
assign weight_0_25[4] = a[4] & b[21];
assign weight_0_25[5] = a[5] & b[20];
assign weight_0_25[6] = a[6] & b[19];
assign weight_0_25[7] = a[7] & b[18];
assign weight_0_25[8] = a[8] & b[17];
assign weight_0_25[9] = a[9] & b[16];
assign weight_0_25[10] = a[10] & b[15];
assign weight_0_25[11] = a[11] & b[14];
assign weight_0_25[12] = a[12] & b[13];
assign weight_0_25[13] = a[13] & b[12];
assign weight_0_25[14] = a[14] & b[11];
assign weight_0_25[15] = a[15] & b[10];
assign weight_0_25[16] = a[16] & b[9];
assign weight_0_25[17] = a[17] & b[8];
assign weight_0_25[18] = a[18] & b[7];
assign weight_0_25[19] = a[19] & b[6];
assign weight_0_25[20] = a[20] & b[5];
assign weight_0_25[21] = a[21] & b[4];
assign weight_0_25[22] = a[22] & b[3];
assign weight_0_25[23] = a[23] & b[2];
assign weight_0_25[24] = a[24] & b[1];
assign weight_0_25[25] = a[25] & b[0];
assign weight_0_26[0] = a[0] & b[26];
assign weight_0_26[1] = a[1] & b[25];
assign weight_0_26[2] = a[2] & b[24];
assign weight_0_26[3] = a[3] & b[23];
assign weight_0_26[4] = a[4] & b[22];
assign weight_0_26[5] = a[5] & b[21];
assign weight_0_26[6] = a[6] & b[20];
assign weight_0_26[7] = a[7] & b[19];
assign weight_0_26[8] = a[8] & b[18];
assign weight_0_26[9] = a[9] & b[17];
assign weight_0_26[10] = a[10] & b[16];
assign weight_0_26[11] = a[11] & b[15];
assign weight_0_26[12] = a[12] & b[14];
assign weight_0_26[13] = a[13] & b[13];
assign weight_0_26[14] = a[14] & b[12];
assign weight_0_26[15] = a[15] & b[11];
assign weight_0_26[16] = a[16] & b[10];
assign weight_0_26[17] = a[17] & b[9];
assign weight_0_26[18] = a[18] & b[8];
assign weight_0_26[19] = a[19] & b[7];
assign weight_0_26[20] = a[20] & b[6];
assign weight_0_26[21] = a[21] & b[5];
assign weight_0_26[22] = a[22] & b[4];
assign weight_0_26[23] = a[23] & b[3];
assign weight_0_26[24] = a[24] & b[2];
assign weight_0_26[25] = a[25] & b[1];
assign weight_0_26[26] = a[26] & b[0];
assign weight_0_27[0] = a[0] & b[27];
assign weight_0_27[1] = a[1] & b[26];
assign weight_0_27[2] = a[2] & b[25];
assign weight_0_27[3] = a[3] & b[24];
assign weight_0_27[4] = a[4] & b[23];
assign weight_0_27[5] = a[5] & b[22];
assign weight_0_27[6] = a[6] & b[21];
assign weight_0_27[7] = a[7] & b[20];
assign weight_0_27[8] = a[8] & b[19];
assign weight_0_27[9] = a[9] & b[18];
assign weight_0_27[10] = a[10] & b[17];
assign weight_0_27[11] = a[11] & b[16];
assign weight_0_27[12] = a[12] & b[15];
assign weight_0_27[13] = a[13] & b[14];
assign weight_0_27[14] = a[14] & b[13];
assign weight_0_27[15] = a[15] & b[12];
assign weight_0_27[16] = a[16] & b[11];
assign weight_0_27[17] = a[17] & b[10];
assign weight_0_27[18] = a[18] & b[9];
assign weight_0_27[19] = a[19] & b[8];
assign weight_0_27[20] = a[20] & b[7];
assign weight_0_27[21] = a[21] & b[6];
assign weight_0_27[22] = a[22] & b[5];
assign weight_0_27[23] = a[23] & b[4];
assign weight_0_27[24] = a[24] & b[3];
assign weight_0_27[25] = a[25] & b[2];
assign weight_0_27[26] = a[26] & b[1];
assign weight_0_27[27] = a[27] & b[0];
assign weight_0_28[0] = a[0] & b[28];
assign weight_0_28[1] = a[1] & b[27];
assign weight_0_28[2] = a[2] & b[26];
assign weight_0_28[3] = a[3] & b[25];
assign weight_0_28[4] = a[4] & b[24];
assign weight_0_28[5] = a[5] & b[23];
assign weight_0_28[6] = a[6] & b[22];
assign weight_0_28[7] = a[7] & b[21];
assign weight_0_28[8] = a[8] & b[20];
assign weight_0_28[9] = a[9] & b[19];
assign weight_0_28[10] = a[10] & b[18];
assign weight_0_28[11] = a[11] & b[17];
assign weight_0_28[12] = a[12] & b[16];
assign weight_0_28[13] = a[13] & b[15];
assign weight_0_28[14] = a[14] & b[14];
assign weight_0_28[15] = a[15] & b[13];
assign weight_0_28[16] = a[16] & b[12];
assign weight_0_28[17] = a[17] & b[11];
assign weight_0_28[18] = a[18] & b[10];
assign weight_0_28[19] = a[19] & b[9];
assign weight_0_28[20] = a[20] & b[8];
assign weight_0_28[21] = a[21] & b[7];
assign weight_0_28[22] = a[22] & b[6];
assign weight_0_28[23] = a[23] & b[5];
assign weight_0_28[24] = a[24] & b[4];
assign weight_0_28[25] = a[25] & b[3];
assign weight_0_28[26] = a[26] & b[2];
assign weight_0_28[27] = a[27] & b[1];
assign weight_0_28[28] = a[28] & b[0];
assign weight_0_29[0] = a[0] & b[29];
assign weight_0_29[1] = a[1] & b[28];
assign weight_0_29[2] = a[2] & b[27];
assign weight_0_29[3] = a[3] & b[26];
assign weight_0_29[4] = a[4] & b[25];
assign weight_0_29[5] = a[5] & b[24];
assign weight_0_29[6] = a[6] & b[23];
assign weight_0_29[7] = a[7] & b[22];
assign weight_0_29[8] = a[8] & b[21];
assign weight_0_29[9] = a[9] & b[20];
assign weight_0_29[10] = a[10] & b[19];
assign weight_0_29[11] = a[11] & b[18];
assign weight_0_29[12] = a[12] & b[17];
assign weight_0_29[13] = a[13] & b[16];
assign weight_0_29[14] = a[14] & b[15];
assign weight_0_29[15] = a[15] & b[14];
assign weight_0_29[16] = a[16] & b[13];
assign weight_0_29[17] = a[17] & b[12];
assign weight_0_29[18] = a[18] & b[11];
assign weight_0_29[19] = a[19] & b[10];
assign weight_0_29[20] = a[20] & b[9];
assign weight_0_29[21] = a[21] & b[8];
assign weight_0_29[22] = a[22] & b[7];
assign weight_0_29[23] = a[23] & b[6];
assign weight_0_29[24] = a[24] & b[5];
assign weight_0_29[25] = a[25] & b[4];
assign weight_0_29[26] = a[26] & b[3];
assign weight_0_29[27] = a[27] & b[2];
assign weight_0_29[28] = a[28] & b[1];
assign weight_0_29[29] = a[29] & b[0];
assign weight_0_30[0] = a[0] & b[30];
assign weight_0_30[1] = a[1] & b[29];
assign weight_0_30[2] = a[2] & b[28];
assign weight_0_30[3] = a[3] & b[27];
assign weight_0_30[4] = a[4] & b[26];
assign weight_0_30[5] = a[5] & b[25];
assign weight_0_30[6] = a[6] & b[24];
assign weight_0_30[7] = a[7] & b[23];
assign weight_0_30[8] = a[8] & b[22];
assign weight_0_30[9] = a[9] & b[21];
assign weight_0_30[10] = a[10] & b[20];
assign weight_0_30[11] = a[11] & b[19];
assign weight_0_30[12] = a[12] & b[18];
assign weight_0_30[13] = a[13] & b[17];
assign weight_0_30[14] = a[14] & b[16];
assign weight_0_30[15] = a[15] & b[15];
assign weight_0_30[16] = a[16] & b[14];
assign weight_0_30[17] = a[17] & b[13];
assign weight_0_30[18] = a[18] & b[12];
assign weight_0_30[19] = a[19] & b[11];
assign weight_0_30[20] = a[20] & b[10];
assign weight_0_30[21] = a[21] & b[9];
assign weight_0_30[22] = a[22] & b[8];
assign weight_0_30[23] = a[23] & b[7];
assign weight_0_30[24] = a[24] & b[6];
assign weight_0_30[25] = a[25] & b[5];
assign weight_0_30[26] = a[26] & b[4];
assign weight_0_30[27] = a[27] & b[3];
assign weight_0_30[28] = a[28] & b[2];
assign weight_0_30[29] = a[29] & b[1];
assign weight_0_30[30] = a[30] & b[0];
assign weight_0_31[0] = a[0] & b[31];
assign weight_0_31[1] = a[1] & b[30];
assign weight_0_31[2] = a[2] & b[29];
assign weight_0_31[3] = a[3] & b[28];
assign weight_0_31[4] = a[4] & b[27];
assign weight_0_31[5] = a[5] & b[26];
assign weight_0_31[6] = a[6] & b[25];
assign weight_0_31[7] = a[7] & b[24];
assign weight_0_31[8] = a[8] & b[23];
assign weight_0_31[9] = a[9] & b[22];
assign weight_0_31[10] = a[10] & b[21];
assign weight_0_31[11] = a[11] & b[20];
assign weight_0_31[12] = a[12] & b[19];
assign weight_0_31[13] = a[13] & b[18];
assign weight_0_31[14] = a[14] & b[17];
assign weight_0_31[15] = a[15] & b[16];
assign weight_0_31[16] = a[16] & b[15];
assign weight_0_31[17] = a[17] & b[14];
assign weight_0_31[18] = a[18] & b[13];
assign weight_0_31[19] = a[19] & b[12];
assign weight_0_31[20] = a[20] & b[11];
assign weight_0_31[21] = a[21] & b[10];
assign weight_0_31[22] = a[22] & b[9];
assign weight_0_31[23] = a[23] & b[8];
assign weight_0_31[24] = a[24] & b[7];
assign weight_0_31[25] = a[25] & b[6];
assign weight_0_31[26] = a[26] & b[5];
assign weight_0_31[27] = a[27] & b[4];
assign weight_0_31[28] = a[28] & b[3];
assign weight_0_31[29] = a[29] & b[2];
assign weight_0_31[30] = a[30] & b[1];
assign weight_0_31[31] = a[31] & b[0];
assign weight_0_32[0] = a[1] & b[31];
assign weight_0_32[1] = a[2] & b[30];
assign weight_0_32[2] = a[3] & b[29];
assign weight_0_32[3] = a[4] & b[28];
assign weight_0_32[4] = a[5] & b[27];
assign weight_0_32[5] = a[6] & b[26];
assign weight_0_32[6] = a[7] & b[25];
assign weight_0_32[7] = a[8] & b[24];
assign weight_0_32[8] = a[9] & b[23];
assign weight_0_32[9] = a[10] & b[22];
assign weight_0_32[10] = a[11] & b[21];
assign weight_0_32[11] = a[12] & b[20];
assign weight_0_32[12] = a[13] & b[19];
assign weight_0_32[13] = a[14] & b[18];
assign weight_0_32[14] = a[15] & b[17];
assign weight_0_32[15] = a[16] & b[16];
assign weight_0_32[16] = a[17] & b[15];
assign weight_0_32[17] = a[18] & b[14];
assign weight_0_32[18] = a[19] & b[13];
assign weight_0_32[19] = a[20] & b[12];
assign weight_0_32[20] = a[21] & b[11];
assign weight_0_32[21] = a[22] & b[10];
assign weight_0_32[22] = a[23] & b[9];
assign weight_0_32[23] = a[24] & b[8];
assign weight_0_32[24] = a[25] & b[7];
assign weight_0_32[25] = a[26] & b[6];
assign weight_0_32[26] = a[27] & b[5];
assign weight_0_32[27] = a[28] & b[4];
assign weight_0_32[28] = a[29] & b[3];
assign weight_0_32[29] = a[30] & b[2];
assign weight_0_32[30] = a[31] & b[1];
assign weight_0_33[0] = a[2] & b[31];
assign weight_0_33[1] = a[3] & b[30];
assign weight_0_33[2] = a[4] & b[29];
assign weight_0_33[3] = a[5] & b[28];
assign weight_0_33[4] = a[6] & b[27];
assign weight_0_33[5] = a[7] & b[26];
assign weight_0_33[6] = a[8] & b[25];
assign weight_0_33[7] = a[9] & b[24];
assign weight_0_33[8] = a[10] & b[23];
assign weight_0_33[9] = a[11] & b[22];
assign weight_0_33[10] = a[12] & b[21];
assign weight_0_33[11] = a[13] & b[20];
assign weight_0_33[12] = a[14] & b[19];
assign weight_0_33[13] = a[15] & b[18];
assign weight_0_33[14] = a[16] & b[17];
assign weight_0_33[15] = a[17] & b[16];
assign weight_0_33[16] = a[18] & b[15];
assign weight_0_33[17] = a[19] & b[14];
assign weight_0_33[18] = a[20] & b[13];
assign weight_0_33[19] = a[21] & b[12];
assign weight_0_33[20] = a[22] & b[11];
assign weight_0_33[21] = a[23] & b[10];
assign weight_0_33[22] = a[24] & b[9];
assign weight_0_33[23] = a[25] & b[8];
assign weight_0_33[24] = a[26] & b[7];
assign weight_0_33[25] = a[27] & b[6];
assign weight_0_33[26] = a[28] & b[5];
assign weight_0_33[27] = a[29] & b[4];
assign weight_0_33[28] = a[30] & b[3];
assign weight_0_33[29] = a[31] & b[2];
assign weight_0_34[0] = a[3] & b[31];
assign weight_0_34[1] = a[4] & b[30];
assign weight_0_34[2] = a[5] & b[29];
assign weight_0_34[3] = a[6] & b[28];
assign weight_0_34[4] = a[7] & b[27];
assign weight_0_34[5] = a[8] & b[26];
assign weight_0_34[6] = a[9] & b[25];
assign weight_0_34[7] = a[10] & b[24];
assign weight_0_34[8] = a[11] & b[23];
assign weight_0_34[9] = a[12] & b[22];
assign weight_0_34[10] = a[13] & b[21];
assign weight_0_34[11] = a[14] & b[20];
assign weight_0_34[12] = a[15] & b[19];
assign weight_0_34[13] = a[16] & b[18];
assign weight_0_34[14] = a[17] & b[17];
assign weight_0_34[15] = a[18] & b[16];
assign weight_0_34[16] = a[19] & b[15];
assign weight_0_34[17] = a[20] & b[14];
assign weight_0_34[18] = a[21] & b[13];
assign weight_0_34[19] = a[22] & b[12];
assign weight_0_34[20] = a[23] & b[11];
assign weight_0_34[21] = a[24] & b[10];
assign weight_0_34[22] = a[25] & b[9];
assign weight_0_34[23] = a[26] & b[8];
assign weight_0_34[24] = a[27] & b[7];
assign weight_0_34[25] = a[28] & b[6];
assign weight_0_34[26] = a[29] & b[5];
assign weight_0_34[27] = a[30] & b[4];
assign weight_0_34[28] = a[31] & b[3];
assign weight_0_35[0] = a[4] & b[31];
assign weight_0_35[1] = a[5] & b[30];
assign weight_0_35[2] = a[6] & b[29];
assign weight_0_35[3] = a[7] & b[28];
assign weight_0_35[4] = a[8] & b[27];
assign weight_0_35[5] = a[9] & b[26];
assign weight_0_35[6] = a[10] & b[25];
assign weight_0_35[7] = a[11] & b[24];
assign weight_0_35[8] = a[12] & b[23];
assign weight_0_35[9] = a[13] & b[22];
assign weight_0_35[10] = a[14] & b[21];
assign weight_0_35[11] = a[15] & b[20];
assign weight_0_35[12] = a[16] & b[19];
assign weight_0_35[13] = a[17] & b[18];
assign weight_0_35[14] = a[18] & b[17];
assign weight_0_35[15] = a[19] & b[16];
assign weight_0_35[16] = a[20] & b[15];
assign weight_0_35[17] = a[21] & b[14];
assign weight_0_35[18] = a[22] & b[13];
assign weight_0_35[19] = a[23] & b[12];
assign weight_0_35[20] = a[24] & b[11];
assign weight_0_35[21] = a[25] & b[10];
assign weight_0_35[22] = a[26] & b[9];
assign weight_0_35[23] = a[27] & b[8];
assign weight_0_35[24] = a[28] & b[7];
assign weight_0_35[25] = a[29] & b[6];
assign weight_0_35[26] = a[30] & b[5];
assign weight_0_35[27] = a[31] & b[4];
assign weight_0_36[0] = a[5] & b[31];
assign weight_0_36[1] = a[6] & b[30];
assign weight_0_36[2] = a[7] & b[29];
assign weight_0_36[3] = a[8] & b[28];
assign weight_0_36[4] = a[9] & b[27];
assign weight_0_36[5] = a[10] & b[26];
assign weight_0_36[6] = a[11] & b[25];
assign weight_0_36[7] = a[12] & b[24];
assign weight_0_36[8] = a[13] & b[23];
assign weight_0_36[9] = a[14] & b[22];
assign weight_0_36[10] = a[15] & b[21];
assign weight_0_36[11] = a[16] & b[20];
assign weight_0_36[12] = a[17] & b[19];
assign weight_0_36[13] = a[18] & b[18];
assign weight_0_36[14] = a[19] & b[17];
assign weight_0_36[15] = a[20] & b[16];
assign weight_0_36[16] = a[21] & b[15];
assign weight_0_36[17] = a[22] & b[14];
assign weight_0_36[18] = a[23] & b[13];
assign weight_0_36[19] = a[24] & b[12];
assign weight_0_36[20] = a[25] & b[11];
assign weight_0_36[21] = a[26] & b[10];
assign weight_0_36[22] = a[27] & b[9];
assign weight_0_36[23] = a[28] & b[8];
assign weight_0_36[24] = a[29] & b[7];
assign weight_0_36[25] = a[30] & b[6];
assign weight_0_36[26] = a[31] & b[5];
assign weight_0_37[0] = a[6] & b[31];
assign weight_0_37[1] = a[7] & b[30];
assign weight_0_37[2] = a[8] & b[29];
assign weight_0_37[3] = a[9] & b[28];
assign weight_0_37[4] = a[10] & b[27];
assign weight_0_37[5] = a[11] & b[26];
assign weight_0_37[6] = a[12] & b[25];
assign weight_0_37[7] = a[13] & b[24];
assign weight_0_37[8] = a[14] & b[23];
assign weight_0_37[9] = a[15] & b[22];
assign weight_0_37[10] = a[16] & b[21];
assign weight_0_37[11] = a[17] & b[20];
assign weight_0_37[12] = a[18] & b[19];
assign weight_0_37[13] = a[19] & b[18];
assign weight_0_37[14] = a[20] & b[17];
assign weight_0_37[15] = a[21] & b[16];
assign weight_0_37[16] = a[22] & b[15];
assign weight_0_37[17] = a[23] & b[14];
assign weight_0_37[18] = a[24] & b[13];
assign weight_0_37[19] = a[25] & b[12];
assign weight_0_37[20] = a[26] & b[11];
assign weight_0_37[21] = a[27] & b[10];
assign weight_0_37[22] = a[28] & b[9];
assign weight_0_37[23] = a[29] & b[8];
assign weight_0_37[24] = a[30] & b[7];
assign weight_0_37[25] = a[31] & b[6];
assign weight_0_38[0] = a[7] & b[31];
assign weight_0_38[1] = a[8] & b[30];
assign weight_0_38[2] = a[9] & b[29];
assign weight_0_38[3] = a[10] & b[28];
assign weight_0_38[4] = a[11] & b[27];
assign weight_0_38[5] = a[12] & b[26];
assign weight_0_38[6] = a[13] & b[25];
assign weight_0_38[7] = a[14] & b[24];
assign weight_0_38[8] = a[15] & b[23];
assign weight_0_38[9] = a[16] & b[22];
assign weight_0_38[10] = a[17] & b[21];
assign weight_0_38[11] = a[18] & b[20];
assign weight_0_38[12] = a[19] & b[19];
assign weight_0_38[13] = a[20] & b[18];
assign weight_0_38[14] = a[21] & b[17];
assign weight_0_38[15] = a[22] & b[16];
assign weight_0_38[16] = a[23] & b[15];
assign weight_0_38[17] = a[24] & b[14];
assign weight_0_38[18] = a[25] & b[13];
assign weight_0_38[19] = a[26] & b[12];
assign weight_0_38[20] = a[27] & b[11];
assign weight_0_38[21] = a[28] & b[10];
assign weight_0_38[22] = a[29] & b[9];
assign weight_0_38[23] = a[30] & b[8];
assign weight_0_38[24] = a[31] & b[7];
assign weight_0_39[0] = a[8] & b[31];
assign weight_0_39[1] = a[9] & b[30];
assign weight_0_39[2] = a[10] & b[29];
assign weight_0_39[3] = a[11] & b[28];
assign weight_0_39[4] = a[12] & b[27];
assign weight_0_39[5] = a[13] & b[26];
assign weight_0_39[6] = a[14] & b[25];
assign weight_0_39[7] = a[15] & b[24];
assign weight_0_39[8] = a[16] & b[23];
assign weight_0_39[9] = a[17] & b[22];
assign weight_0_39[10] = a[18] & b[21];
assign weight_0_39[11] = a[19] & b[20];
assign weight_0_39[12] = a[20] & b[19];
assign weight_0_39[13] = a[21] & b[18];
assign weight_0_39[14] = a[22] & b[17];
assign weight_0_39[15] = a[23] & b[16];
assign weight_0_39[16] = a[24] & b[15];
assign weight_0_39[17] = a[25] & b[14];
assign weight_0_39[18] = a[26] & b[13];
assign weight_0_39[19] = a[27] & b[12];
assign weight_0_39[20] = a[28] & b[11];
assign weight_0_39[21] = a[29] & b[10];
assign weight_0_39[22] = a[30] & b[9];
assign weight_0_39[23] = a[31] & b[8];
assign weight_0_40[0] = a[9] & b[31];
assign weight_0_40[1] = a[10] & b[30];
assign weight_0_40[2] = a[11] & b[29];
assign weight_0_40[3] = a[12] & b[28];
assign weight_0_40[4] = a[13] & b[27];
assign weight_0_40[5] = a[14] & b[26];
assign weight_0_40[6] = a[15] & b[25];
assign weight_0_40[7] = a[16] & b[24];
assign weight_0_40[8] = a[17] & b[23];
assign weight_0_40[9] = a[18] & b[22];
assign weight_0_40[10] = a[19] & b[21];
assign weight_0_40[11] = a[20] & b[20];
assign weight_0_40[12] = a[21] & b[19];
assign weight_0_40[13] = a[22] & b[18];
assign weight_0_40[14] = a[23] & b[17];
assign weight_0_40[15] = a[24] & b[16];
assign weight_0_40[16] = a[25] & b[15];
assign weight_0_40[17] = a[26] & b[14];
assign weight_0_40[18] = a[27] & b[13];
assign weight_0_40[19] = a[28] & b[12];
assign weight_0_40[20] = a[29] & b[11];
assign weight_0_40[21] = a[30] & b[10];
assign weight_0_40[22] = a[31] & b[9];
assign weight_0_41[0] = a[10] & b[31];
assign weight_0_41[1] = a[11] & b[30];
assign weight_0_41[2] = a[12] & b[29];
assign weight_0_41[3] = a[13] & b[28];
assign weight_0_41[4] = a[14] & b[27];
assign weight_0_41[5] = a[15] & b[26];
assign weight_0_41[6] = a[16] & b[25];
assign weight_0_41[7] = a[17] & b[24];
assign weight_0_41[8] = a[18] & b[23];
assign weight_0_41[9] = a[19] & b[22];
assign weight_0_41[10] = a[20] & b[21];
assign weight_0_41[11] = a[21] & b[20];
assign weight_0_41[12] = a[22] & b[19];
assign weight_0_41[13] = a[23] & b[18];
assign weight_0_41[14] = a[24] & b[17];
assign weight_0_41[15] = a[25] & b[16];
assign weight_0_41[16] = a[26] & b[15];
assign weight_0_41[17] = a[27] & b[14];
assign weight_0_41[18] = a[28] & b[13];
assign weight_0_41[19] = a[29] & b[12];
assign weight_0_41[20] = a[30] & b[11];
assign weight_0_41[21] = a[31] & b[10];
assign weight_0_42[0] = a[11] & b[31];
assign weight_0_42[1] = a[12] & b[30];
assign weight_0_42[2] = a[13] & b[29];
assign weight_0_42[3] = a[14] & b[28];
assign weight_0_42[4] = a[15] & b[27];
assign weight_0_42[5] = a[16] & b[26];
assign weight_0_42[6] = a[17] & b[25];
assign weight_0_42[7] = a[18] & b[24];
assign weight_0_42[8] = a[19] & b[23];
assign weight_0_42[9] = a[20] & b[22];
assign weight_0_42[10] = a[21] & b[21];
assign weight_0_42[11] = a[22] & b[20];
assign weight_0_42[12] = a[23] & b[19];
assign weight_0_42[13] = a[24] & b[18];
assign weight_0_42[14] = a[25] & b[17];
assign weight_0_42[15] = a[26] & b[16];
assign weight_0_42[16] = a[27] & b[15];
assign weight_0_42[17] = a[28] & b[14];
assign weight_0_42[18] = a[29] & b[13];
assign weight_0_42[19] = a[30] & b[12];
assign weight_0_42[20] = a[31] & b[11];
assign weight_0_43[0] = a[12] & b[31];
assign weight_0_43[1] = a[13] & b[30];
assign weight_0_43[2] = a[14] & b[29];
assign weight_0_43[3] = a[15] & b[28];
assign weight_0_43[4] = a[16] & b[27];
assign weight_0_43[5] = a[17] & b[26];
assign weight_0_43[6] = a[18] & b[25];
assign weight_0_43[7] = a[19] & b[24];
assign weight_0_43[8] = a[20] & b[23];
assign weight_0_43[9] = a[21] & b[22];
assign weight_0_43[10] = a[22] & b[21];
assign weight_0_43[11] = a[23] & b[20];
assign weight_0_43[12] = a[24] & b[19];
assign weight_0_43[13] = a[25] & b[18];
assign weight_0_43[14] = a[26] & b[17];
assign weight_0_43[15] = a[27] & b[16];
assign weight_0_43[16] = a[28] & b[15];
assign weight_0_43[17] = a[29] & b[14];
assign weight_0_43[18] = a[30] & b[13];
assign weight_0_43[19] = a[31] & b[12];
assign weight_0_44[0] = a[13] & b[31];
assign weight_0_44[1] = a[14] & b[30];
assign weight_0_44[2] = a[15] & b[29];
assign weight_0_44[3] = a[16] & b[28];
assign weight_0_44[4] = a[17] & b[27];
assign weight_0_44[5] = a[18] & b[26];
assign weight_0_44[6] = a[19] & b[25];
assign weight_0_44[7] = a[20] & b[24];
assign weight_0_44[8] = a[21] & b[23];
assign weight_0_44[9] = a[22] & b[22];
assign weight_0_44[10] = a[23] & b[21];
assign weight_0_44[11] = a[24] & b[20];
assign weight_0_44[12] = a[25] & b[19];
assign weight_0_44[13] = a[26] & b[18];
assign weight_0_44[14] = a[27] & b[17];
assign weight_0_44[15] = a[28] & b[16];
assign weight_0_44[16] = a[29] & b[15];
assign weight_0_44[17] = a[30] & b[14];
assign weight_0_44[18] = a[31] & b[13];
assign weight_0_45[0] = a[14] & b[31];
assign weight_0_45[1] = a[15] & b[30];
assign weight_0_45[2] = a[16] & b[29];
assign weight_0_45[3] = a[17] & b[28];
assign weight_0_45[4] = a[18] & b[27];
assign weight_0_45[5] = a[19] & b[26];
assign weight_0_45[6] = a[20] & b[25];
assign weight_0_45[7] = a[21] & b[24];
assign weight_0_45[8] = a[22] & b[23];
assign weight_0_45[9] = a[23] & b[22];
assign weight_0_45[10] = a[24] & b[21];
assign weight_0_45[11] = a[25] & b[20];
assign weight_0_45[12] = a[26] & b[19];
assign weight_0_45[13] = a[27] & b[18];
assign weight_0_45[14] = a[28] & b[17];
assign weight_0_45[15] = a[29] & b[16];
assign weight_0_45[16] = a[30] & b[15];
assign weight_0_45[17] = a[31] & b[14];
assign weight_0_46[0] = a[15] & b[31];
assign weight_0_46[1] = a[16] & b[30];
assign weight_0_46[2] = a[17] & b[29];
assign weight_0_46[3] = a[18] & b[28];
assign weight_0_46[4] = a[19] & b[27];
assign weight_0_46[5] = a[20] & b[26];
assign weight_0_46[6] = a[21] & b[25];
assign weight_0_46[7] = a[22] & b[24];
assign weight_0_46[8] = a[23] & b[23];
assign weight_0_46[9] = a[24] & b[22];
assign weight_0_46[10] = a[25] & b[21];
assign weight_0_46[11] = a[26] & b[20];
assign weight_0_46[12] = a[27] & b[19];
assign weight_0_46[13] = a[28] & b[18];
assign weight_0_46[14] = a[29] & b[17];
assign weight_0_46[15] = a[30] & b[16];
assign weight_0_46[16] = a[31] & b[15];
assign weight_0_47[0] = a[16] & b[31];
assign weight_0_47[1] = a[17] & b[30];
assign weight_0_47[2] = a[18] & b[29];
assign weight_0_47[3] = a[19] & b[28];
assign weight_0_47[4] = a[20] & b[27];
assign weight_0_47[5] = a[21] & b[26];
assign weight_0_47[6] = a[22] & b[25];
assign weight_0_47[7] = a[23] & b[24];
assign weight_0_47[8] = a[24] & b[23];
assign weight_0_47[9] = a[25] & b[22];
assign weight_0_47[10] = a[26] & b[21];
assign weight_0_47[11] = a[27] & b[20];
assign weight_0_47[12] = a[28] & b[19];
assign weight_0_47[13] = a[29] & b[18];
assign weight_0_47[14] = a[30] & b[17];
assign weight_0_47[15] = a[31] & b[16];
assign weight_0_48[0] = a[17] & b[31];
assign weight_0_48[1] = a[18] & b[30];
assign weight_0_48[2] = a[19] & b[29];
assign weight_0_48[3] = a[20] & b[28];
assign weight_0_48[4] = a[21] & b[27];
assign weight_0_48[5] = a[22] & b[26];
assign weight_0_48[6] = a[23] & b[25];
assign weight_0_48[7] = a[24] & b[24];
assign weight_0_48[8] = a[25] & b[23];
assign weight_0_48[9] = a[26] & b[22];
assign weight_0_48[10] = a[27] & b[21];
assign weight_0_48[11] = a[28] & b[20];
assign weight_0_48[12] = a[29] & b[19];
assign weight_0_48[13] = a[30] & b[18];
assign weight_0_48[14] = a[31] & b[17];
assign weight_0_49[0] = a[18] & b[31];
assign weight_0_49[1] = a[19] & b[30];
assign weight_0_49[2] = a[20] & b[29];
assign weight_0_49[3] = a[21] & b[28];
assign weight_0_49[4] = a[22] & b[27];
assign weight_0_49[5] = a[23] & b[26];
assign weight_0_49[6] = a[24] & b[25];
assign weight_0_49[7] = a[25] & b[24];
assign weight_0_49[8] = a[26] & b[23];
assign weight_0_49[9] = a[27] & b[22];
assign weight_0_49[10] = a[28] & b[21];
assign weight_0_49[11] = a[29] & b[20];
assign weight_0_49[12] = a[30] & b[19];
assign weight_0_49[13] = a[31] & b[18];
assign weight_0_50[0] = a[19] & b[31];
assign weight_0_50[1] = a[20] & b[30];
assign weight_0_50[2] = a[21] & b[29];
assign weight_0_50[3] = a[22] & b[28];
assign weight_0_50[4] = a[23] & b[27];
assign weight_0_50[5] = a[24] & b[26];
assign weight_0_50[6] = a[25] & b[25];
assign weight_0_50[7] = a[26] & b[24];
assign weight_0_50[8] = a[27] & b[23];
assign weight_0_50[9] = a[28] & b[22];
assign weight_0_50[10] = a[29] & b[21];
assign weight_0_50[11] = a[30] & b[20];
assign weight_0_50[12] = a[31] & b[19];
assign weight_0_51[0] = a[20] & b[31];
assign weight_0_51[1] = a[21] & b[30];
assign weight_0_51[2] = a[22] & b[29];
assign weight_0_51[3] = a[23] & b[28];
assign weight_0_51[4] = a[24] & b[27];
assign weight_0_51[5] = a[25] & b[26];
assign weight_0_51[6] = a[26] & b[25];
assign weight_0_51[7] = a[27] & b[24];
assign weight_0_51[8] = a[28] & b[23];
assign weight_0_51[9] = a[29] & b[22];
assign weight_0_51[10] = a[30] & b[21];
assign weight_0_51[11] = a[31] & b[20];
assign weight_0_52[0] = a[21] & b[31];
assign weight_0_52[1] = a[22] & b[30];
assign weight_0_52[2] = a[23] & b[29];
assign weight_0_52[3] = a[24] & b[28];
assign weight_0_52[4] = a[25] & b[27];
assign weight_0_52[5] = a[26] & b[26];
assign weight_0_52[6] = a[27] & b[25];
assign weight_0_52[7] = a[28] & b[24];
assign weight_0_52[8] = a[29] & b[23];
assign weight_0_52[9] = a[30] & b[22];
assign weight_0_52[10] = a[31] & b[21];
assign weight_0_53[0] = a[22] & b[31];
assign weight_0_53[1] = a[23] & b[30];
assign weight_0_53[2] = a[24] & b[29];
assign weight_0_53[3] = a[25] & b[28];
assign weight_0_53[4] = a[26] & b[27];
assign weight_0_53[5] = a[27] & b[26];
assign weight_0_53[6] = a[28] & b[25];
assign weight_0_53[7] = a[29] & b[24];
assign weight_0_53[8] = a[30] & b[23];
assign weight_0_53[9] = a[31] & b[22];
assign weight_0_54[0] = a[23] & b[31];
assign weight_0_54[1] = a[24] & b[30];
assign weight_0_54[2] = a[25] & b[29];
assign weight_0_54[3] = a[26] & b[28];
assign weight_0_54[4] = a[27] & b[27];
assign weight_0_54[5] = a[28] & b[26];
assign weight_0_54[6] = a[29] & b[25];
assign weight_0_54[7] = a[30] & b[24];
assign weight_0_54[8] = a[31] & b[23];
assign weight_0_55[0] = a[24] & b[31];
assign weight_0_55[1] = a[25] & b[30];
assign weight_0_55[2] = a[26] & b[29];
assign weight_0_55[3] = a[27] & b[28];
assign weight_0_55[4] = a[28] & b[27];
assign weight_0_55[5] = a[29] & b[26];
assign weight_0_55[6] = a[30] & b[25];
assign weight_0_55[7] = a[31] & b[24];
assign weight_0_56[0] = a[25] & b[31];
assign weight_0_56[1] = a[26] & b[30];
assign weight_0_56[2] = a[27] & b[29];
assign weight_0_56[3] = a[28] & b[28];
assign weight_0_56[4] = a[29] & b[27];
assign weight_0_56[5] = a[30] & b[26];
assign weight_0_56[6] = a[31] & b[25];
assign weight_0_57[0] = a[26] & b[31];
assign weight_0_57[1] = a[27] & b[30];
assign weight_0_57[2] = a[28] & b[29];
assign weight_0_57[3] = a[29] & b[28];
assign weight_0_57[4] = a[30] & b[27];
assign weight_0_57[5] = a[31] & b[26];
assign weight_0_58[0] = a[27] & b[31];
assign weight_0_58[1] = a[28] & b[30];
assign weight_0_58[2] = a[29] & b[29];
assign weight_0_58[3] = a[30] & b[28];
assign weight_0_58[4] = a[31] & b[27];
assign weight_0_59[0] = a[28] & b[31];
assign weight_0_59[1] = a[29] & b[30];
assign weight_0_59[2] = a[30] & b[29];
assign weight_0_59[3] = a[31] & b[28];
assign weight_0_60[0] = a[29] & b[31];
assign weight_0_60[1] = a[30] & b[30];
assign weight_0_60[2] = a[31] & b[29];
assign weight_0_61[0] = a[30] & b[31];
assign weight_0_61[1] = a[31] & b[30];
assign weight_0_62 = a[31] & b[31];
logic weight_1_0;
logic weight_1_1;
logic [1:0] weight_1_2;
logic [2:0] weight_1_3;
logic [2:0] weight_1_4;
logic [3:0] weight_1_5;
logic [4:0] weight_1_6;
logic [4:0] weight_1_7;
logic [5:0] weight_1_8;
logic [6:0] weight_1_9;
logic [6:0] weight_1_10;
logic [7:0] weight_1_11;
logic [8:0] weight_1_12;
logic [8:0] weight_1_13;
logic [9:0] weight_1_14;
logic [10:0] weight_1_15;
logic [10:0] weight_1_16;
logic [11:0] weight_1_17;
logic [12:0] weight_1_18;
logic [12:0] weight_1_19;
logic [13:0] weight_1_20;
logic [14:0] weight_1_21;
logic [14:0] weight_1_22;
logic [15:0] weight_1_23;
logic [16:0] weight_1_24;
logic [16:0] weight_1_25;
logic [17:0] weight_1_26;
logic [18:0] weight_1_27;
logic [18:0] weight_1_28;
logic [19:0] weight_1_29;
logic [20:0] weight_1_30;
logic [21:0] weight_1_31;
logic [21:0] weight_1_32;
logic [21:0] weight_1_33;
logic [19:0] weight_1_34;
logic [19:0] weight_1_35;
logic [19:0] weight_1_36;
logic [17:0] weight_1_37;
logic [17:0] weight_1_38;
logic [17:0] weight_1_39;
logic [15:0] weight_1_40;
logic [15:0] weight_1_41;
logic [15:0] weight_1_42;
logic [13:0] weight_1_43;
logic [13:0] weight_1_44;
logic [13:0] weight_1_45;
logic [11:0] weight_1_46;
logic [11:0] weight_1_47;
logic [11:0] weight_1_48;
logic [9:0] weight_1_49;
logic [9:0] weight_1_50;
logic [9:0] weight_1_51;
logic [7:0] weight_1_52;
logic [7:0] weight_1_53;
logic [7:0] weight_1_54;
logic [5:0] weight_1_55;
logic [5:0] weight_1_56;
logic [5:0] weight_1_57;
logic [3:0] weight_1_58;
logic [3:0] weight_1_59;
logic [3:0] weight_1_60;
logic [1:0] weight_1_61;
logic weight_1_62;
assign weight_1_0 = weight_0_0;
half_adder ha0(.a(weight_0_1[0]), .b(weight_0_1[1]), .sum(weight_1_1), .cout(weight_1_2[0]));
full_adder fa0(.a(weight_0_2[0]), .b(weight_0_2[1]), .cin(weight_0_2[2]), .sum(weight_1_2[1]), .cout(weight_1_3[0]));
full_adder fa1(.a(weight_0_3[0]), .b(weight_0_3[1]), .cin(weight_0_3[2]), .sum(weight_1_3[1]), .cout(weight_1_4[0]));
full_adder fa2(.a(weight_0_4[0]), .b(weight_0_4[1]), .cin(weight_0_4[2]), .sum(weight_1_4[1]), .cout(weight_1_5[0]));
full_adder fa3(.a(weight_0_5[0]), .b(weight_0_5[1]), .cin(weight_0_5[2]), .sum(weight_1_5[1]), .cout(weight_1_6[0]));
full_adder fa4(.a(weight_0_6[0]), .b(weight_0_6[1]), .cin(weight_0_6[2]), .sum(weight_1_6[1]), .cout(weight_1_7[0]));
full_adder fa5(.a(weight_0_7[0]), .b(weight_0_7[1]), .cin(weight_0_7[2]), .sum(weight_1_7[1]), .cout(weight_1_8[0]));
full_adder fa6(.a(weight_0_8[0]), .b(weight_0_8[1]), .cin(weight_0_8[2]), .sum(weight_1_8[1]), .cout(weight_1_9[0]));
full_adder fa7(.a(weight_0_9[0]), .b(weight_0_9[1]), .cin(weight_0_9[2]), .sum(weight_1_9[1]), .cout(weight_1_10[0]));
full_adder fa8(.a(weight_0_10[0]), .b(weight_0_10[1]), .cin(weight_0_10[2]), .sum(weight_1_10[1]), .cout(weight_1_11[0]));
full_adder fa9(.a(weight_0_11[0]), .b(weight_0_11[1]), .cin(weight_0_11[2]), .sum(weight_1_11[1]), .cout(weight_1_12[0]));
full_adder fa10(.a(weight_0_12[0]), .b(weight_0_12[1]), .cin(weight_0_12[2]), .sum(weight_1_12[1]), .cout(weight_1_13[0]));
full_adder fa11(.a(weight_0_13[0]), .b(weight_0_13[1]), .cin(weight_0_13[2]), .sum(weight_1_13[1]), .cout(weight_1_14[0]));
full_adder fa12(.a(weight_0_14[0]), .b(weight_0_14[1]), .cin(weight_0_14[2]), .sum(weight_1_14[1]), .cout(weight_1_15[0]));
full_adder fa13(.a(weight_0_15[0]), .b(weight_0_15[1]), .cin(weight_0_15[2]), .sum(weight_1_15[1]), .cout(weight_1_16[0]));
full_adder fa14(.a(weight_0_16[0]), .b(weight_0_16[1]), .cin(weight_0_16[2]), .sum(weight_1_16[1]), .cout(weight_1_17[0]));
full_adder fa15(.a(weight_0_17[0]), .b(weight_0_17[1]), .cin(weight_0_17[2]), .sum(weight_1_17[1]), .cout(weight_1_18[0]));
full_adder fa16(.a(weight_0_18[0]), .b(weight_0_18[1]), .cin(weight_0_18[2]), .sum(weight_1_18[1]), .cout(weight_1_19[0]));
full_adder fa17(.a(weight_0_19[0]), .b(weight_0_19[1]), .cin(weight_0_19[2]), .sum(weight_1_19[1]), .cout(weight_1_20[0]));
full_adder fa18(.a(weight_0_20[0]), .b(weight_0_20[1]), .cin(weight_0_20[2]), .sum(weight_1_20[1]), .cout(weight_1_21[0]));
full_adder fa19(.a(weight_0_21[0]), .b(weight_0_21[1]), .cin(weight_0_21[2]), .sum(weight_1_21[1]), .cout(weight_1_22[0]));
full_adder fa20(.a(weight_0_22[0]), .b(weight_0_22[1]), .cin(weight_0_22[2]), .sum(weight_1_22[1]), .cout(weight_1_23[0]));
full_adder fa21(.a(weight_0_23[0]), .b(weight_0_23[1]), .cin(weight_0_23[2]), .sum(weight_1_23[1]), .cout(weight_1_24[0]));
full_adder fa22(.a(weight_0_24[0]), .b(weight_0_24[1]), .cin(weight_0_24[2]), .sum(weight_1_24[1]), .cout(weight_1_25[0]));
full_adder fa23(.a(weight_0_25[0]), .b(weight_0_25[1]), .cin(weight_0_25[2]), .sum(weight_1_25[1]), .cout(weight_1_26[0]));
full_adder fa24(.a(weight_0_26[0]), .b(weight_0_26[1]), .cin(weight_0_26[2]), .sum(weight_1_26[1]), .cout(weight_1_27[0]));
full_adder fa25(.a(weight_0_27[0]), .b(weight_0_27[1]), .cin(weight_0_27[2]), .sum(weight_1_27[1]), .cout(weight_1_28[0]));
full_adder fa26(.a(weight_0_28[0]), .b(weight_0_28[1]), .cin(weight_0_28[2]), .sum(weight_1_28[1]), .cout(weight_1_29[0]));
full_adder fa27(.a(weight_0_29[0]), .b(weight_0_29[1]), .cin(weight_0_29[2]), .sum(weight_1_29[1]), .cout(weight_1_30[0]));
full_adder fa28(.a(weight_0_30[0]), .b(weight_0_30[1]), .cin(weight_0_30[2]), .sum(weight_1_30[1]), .cout(weight_1_31[0]));
full_adder fa29(.a(weight_0_31[0]), .b(weight_0_31[1]), .cin(weight_0_31[2]), .sum(weight_1_31[1]), .cout(weight_1_32[0]));
half_adder ha1(.a(weight_0_32[0]), .b(weight_0_32[1]), .sum(weight_1_32[1]), .cout(weight_1_33[0]));
assign weight_1_33[1] = weight_0_33[0];
assign weight_1_3[2] = weight_0_3[3];
half_adder ha2(.a(weight_0_4[3]), .b(weight_0_4[4]), .sum(weight_1_4[2]), .cout(weight_1_5[2]));
full_adder fa30(.a(weight_0_5[3]), .b(weight_0_5[4]), .cin(weight_0_5[5]), .sum(weight_1_5[3]), .cout(weight_1_6[2]));
full_adder fa31(.a(weight_0_6[3]), .b(weight_0_6[4]), .cin(weight_0_6[5]), .sum(weight_1_6[3]), .cout(weight_1_7[2]));
full_adder fa32(.a(weight_0_7[3]), .b(weight_0_7[4]), .cin(weight_0_7[5]), .sum(weight_1_7[3]), .cout(weight_1_8[2]));
full_adder fa33(.a(weight_0_8[3]), .b(weight_0_8[4]), .cin(weight_0_8[5]), .sum(weight_1_8[3]), .cout(weight_1_9[2]));
full_adder fa34(.a(weight_0_9[3]), .b(weight_0_9[4]), .cin(weight_0_9[5]), .sum(weight_1_9[3]), .cout(weight_1_10[2]));
full_adder fa35(.a(weight_0_10[3]), .b(weight_0_10[4]), .cin(weight_0_10[5]), .sum(weight_1_10[3]), .cout(weight_1_11[2]));
full_adder fa36(.a(weight_0_11[3]), .b(weight_0_11[4]), .cin(weight_0_11[5]), .sum(weight_1_11[3]), .cout(weight_1_12[2]));
full_adder fa37(.a(weight_0_12[3]), .b(weight_0_12[4]), .cin(weight_0_12[5]), .sum(weight_1_12[3]), .cout(weight_1_13[2]));
full_adder fa38(.a(weight_0_13[3]), .b(weight_0_13[4]), .cin(weight_0_13[5]), .sum(weight_1_13[3]), .cout(weight_1_14[2]));
full_adder fa39(.a(weight_0_14[3]), .b(weight_0_14[4]), .cin(weight_0_14[5]), .sum(weight_1_14[3]), .cout(weight_1_15[2]));
full_adder fa40(.a(weight_0_15[3]), .b(weight_0_15[4]), .cin(weight_0_15[5]), .sum(weight_1_15[3]), .cout(weight_1_16[2]));
full_adder fa41(.a(weight_0_16[3]), .b(weight_0_16[4]), .cin(weight_0_16[5]), .sum(weight_1_16[3]), .cout(weight_1_17[2]));
full_adder fa42(.a(weight_0_17[3]), .b(weight_0_17[4]), .cin(weight_0_17[5]), .sum(weight_1_17[3]), .cout(weight_1_18[2]));
full_adder fa43(.a(weight_0_18[3]), .b(weight_0_18[4]), .cin(weight_0_18[5]), .sum(weight_1_18[3]), .cout(weight_1_19[2]));
full_adder fa44(.a(weight_0_19[3]), .b(weight_0_19[4]), .cin(weight_0_19[5]), .sum(weight_1_19[3]), .cout(weight_1_20[2]));
full_adder fa45(.a(weight_0_20[3]), .b(weight_0_20[4]), .cin(weight_0_20[5]), .sum(weight_1_20[3]), .cout(weight_1_21[2]));
full_adder fa46(.a(weight_0_21[3]), .b(weight_0_21[4]), .cin(weight_0_21[5]), .sum(weight_1_21[3]), .cout(weight_1_22[2]));
full_adder fa47(.a(weight_0_22[3]), .b(weight_0_22[4]), .cin(weight_0_22[5]), .sum(weight_1_22[3]), .cout(weight_1_23[2]));
full_adder fa48(.a(weight_0_23[3]), .b(weight_0_23[4]), .cin(weight_0_23[5]), .sum(weight_1_23[3]), .cout(weight_1_24[2]));
full_adder fa49(.a(weight_0_24[3]), .b(weight_0_24[4]), .cin(weight_0_24[5]), .sum(weight_1_24[3]), .cout(weight_1_25[2]));
full_adder fa50(.a(weight_0_25[3]), .b(weight_0_25[4]), .cin(weight_0_25[5]), .sum(weight_1_25[3]), .cout(weight_1_26[2]));
full_adder fa51(.a(weight_0_26[3]), .b(weight_0_26[4]), .cin(weight_0_26[5]), .sum(weight_1_26[3]), .cout(weight_1_27[2]));
full_adder fa52(.a(weight_0_27[3]), .b(weight_0_27[4]), .cin(weight_0_27[5]), .sum(weight_1_27[3]), .cout(weight_1_28[2]));
full_adder fa53(.a(weight_0_28[3]), .b(weight_0_28[4]), .cin(weight_0_28[5]), .sum(weight_1_28[3]), .cout(weight_1_29[2]));
full_adder fa54(.a(weight_0_29[3]), .b(weight_0_29[4]), .cin(weight_0_29[5]), .sum(weight_1_29[3]), .cout(weight_1_30[2]));
full_adder fa55(.a(weight_0_30[3]), .b(weight_0_30[4]), .cin(weight_0_30[5]), .sum(weight_1_30[3]), .cout(weight_1_31[2]));
full_adder fa56(.a(weight_0_31[3]), .b(weight_0_31[4]), .cin(weight_0_31[5]), .sum(weight_1_31[3]), .cout(weight_1_32[2]));
full_adder fa57(.a(weight_0_32[2]), .b(weight_0_32[3]), .cin(weight_0_32[4]), .sum(weight_1_32[3]), .cout(weight_1_33[2]));
full_adder fa58(.a(weight_0_33[1]), .b(weight_0_33[2]), .cin(weight_0_33[3]), .sum(weight_1_33[3]), .cout(weight_1_34[0]));
full_adder fa59(.a(weight_0_34[0]), .b(weight_0_34[1]), .cin(weight_0_34[2]), .sum(weight_1_34[1]), .cout(weight_1_35[0]));
half_adder ha3(.a(weight_0_35[0]), .b(weight_0_35[1]), .sum(weight_1_35[1]), .cout(weight_1_36[0]));
assign weight_1_36[1] = weight_0_36[0];
assign weight_1_6[4] = weight_0_6[6];
half_adder ha4(.a(weight_0_7[6]), .b(weight_0_7[7]), .sum(weight_1_7[4]), .cout(weight_1_8[4]));
full_adder fa60(.a(weight_0_8[6]), .b(weight_0_8[7]), .cin(weight_0_8[8]), .sum(weight_1_8[5]), .cout(weight_1_9[4]));
full_adder fa61(.a(weight_0_9[6]), .b(weight_0_9[7]), .cin(weight_0_9[8]), .sum(weight_1_9[5]), .cout(weight_1_10[4]));
full_adder fa62(.a(weight_0_10[6]), .b(weight_0_10[7]), .cin(weight_0_10[8]), .sum(weight_1_10[5]), .cout(weight_1_11[4]));
full_adder fa63(.a(weight_0_11[6]), .b(weight_0_11[7]), .cin(weight_0_11[8]), .sum(weight_1_11[5]), .cout(weight_1_12[4]));
full_adder fa64(.a(weight_0_12[6]), .b(weight_0_12[7]), .cin(weight_0_12[8]), .sum(weight_1_12[5]), .cout(weight_1_13[4]));
full_adder fa65(.a(weight_0_13[6]), .b(weight_0_13[7]), .cin(weight_0_13[8]), .sum(weight_1_13[5]), .cout(weight_1_14[4]));
full_adder fa66(.a(weight_0_14[6]), .b(weight_0_14[7]), .cin(weight_0_14[8]), .sum(weight_1_14[5]), .cout(weight_1_15[4]));
full_adder fa67(.a(weight_0_15[6]), .b(weight_0_15[7]), .cin(weight_0_15[8]), .sum(weight_1_15[5]), .cout(weight_1_16[4]));
full_adder fa68(.a(weight_0_16[6]), .b(weight_0_16[7]), .cin(weight_0_16[8]), .sum(weight_1_16[5]), .cout(weight_1_17[4]));
full_adder fa69(.a(weight_0_17[6]), .b(weight_0_17[7]), .cin(weight_0_17[8]), .sum(weight_1_17[5]), .cout(weight_1_18[4]));
full_adder fa70(.a(weight_0_18[6]), .b(weight_0_18[7]), .cin(weight_0_18[8]), .sum(weight_1_18[5]), .cout(weight_1_19[4]));
full_adder fa71(.a(weight_0_19[6]), .b(weight_0_19[7]), .cin(weight_0_19[8]), .sum(weight_1_19[5]), .cout(weight_1_20[4]));
full_adder fa72(.a(weight_0_20[6]), .b(weight_0_20[7]), .cin(weight_0_20[8]), .sum(weight_1_20[5]), .cout(weight_1_21[4]));
full_adder fa73(.a(weight_0_21[6]), .b(weight_0_21[7]), .cin(weight_0_21[8]), .sum(weight_1_21[5]), .cout(weight_1_22[4]));
full_adder fa74(.a(weight_0_22[6]), .b(weight_0_22[7]), .cin(weight_0_22[8]), .sum(weight_1_22[5]), .cout(weight_1_23[4]));
full_adder fa75(.a(weight_0_23[6]), .b(weight_0_23[7]), .cin(weight_0_23[8]), .sum(weight_1_23[5]), .cout(weight_1_24[4]));
full_adder fa76(.a(weight_0_24[6]), .b(weight_0_24[7]), .cin(weight_0_24[8]), .sum(weight_1_24[5]), .cout(weight_1_25[4]));
full_adder fa77(.a(weight_0_25[6]), .b(weight_0_25[7]), .cin(weight_0_25[8]), .sum(weight_1_25[5]), .cout(weight_1_26[4]));
full_adder fa78(.a(weight_0_26[6]), .b(weight_0_26[7]), .cin(weight_0_26[8]), .sum(weight_1_26[5]), .cout(weight_1_27[4]));
full_adder fa79(.a(weight_0_27[6]), .b(weight_0_27[7]), .cin(weight_0_27[8]), .sum(weight_1_27[5]), .cout(weight_1_28[4]));
full_adder fa80(.a(weight_0_28[6]), .b(weight_0_28[7]), .cin(weight_0_28[8]), .sum(weight_1_28[5]), .cout(weight_1_29[4]));
full_adder fa81(.a(weight_0_29[6]), .b(weight_0_29[7]), .cin(weight_0_29[8]), .sum(weight_1_29[5]), .cout(weight_1_30[4]));
full_adder fa82(.a(weight_0_30[6]), .b(weight_0_30[7]), .cin(weight_0_30[8]), .sum(weight_1_30[5]), .cout(weight_1_31[4]));
full_adder fa83(.a(weight_0_31[6]), .b(weight_0_31[7]), .cin(weight_0_31[8]), .sum(weight_1_31[5]), .cout(weight_1_32[4]));
full_adder fa84(.a(weight_0_32[5]), .b(weight_0_32[6]), .cin(weight_0_32[7]), .sum(weight_1_32[5]), .cout(weight_1_33[4]));
full_adder fa85(.a(weight_0_33[4]), .b(weight_0_33[5]), .cin(weight_0_33[6]), .sum(weight_1_33[5]), .cout(weight_1_34[2]));
full_adder fa86(.a(weight_0_34[3]), .b(weight_0_34[4]), .cin(weight_0_34[5]), .sum(weight_1_34[3]), .cout(weight_1_35[2]));
full_adder fa87(.a(weight_0_35[2]), .b(weight_0_35[3]), .cin(weight_0_35[4]), .sum(weight_1_35[3]), .cout(weight_1_36[2]));
full_adder fa88(.a(weight_0_36[1]), .b(weight_0_36[2]), .cin(weight_0_36[3]), .sum(weight_1_36[3]), .cout(weight_1_37[0]));
full_adder fa89(.a(weight_0_37[0]), .b(weight_0_37[1]), .cin(weight_0_37[2]), .sum(weight_1_37[1]), .cout(weight_1_38[0]));
half_adder ha5(.a(weight_0_38[0]), .b(weight_0_38[1]), .sum(weight_1_38[1]), .cout(weight_1_39[0]));
assign weight_1_39[1] = weight_0_39[0];
assign weight_1_9[6] = weight_0_9[9];
half_adder ha6(.a(weight_0_10[9]), .b(weight_0_10[10]), .sum(weight_1_10[6]), .cout(weight_1_11[6]));
full_adder fa90(.a(weight_0_11[9]), .b(weight_0_11[10]), .cin(weight_0_11[11]), .sum(weight_1_11[7]), .cout(weight_1_12[6]));
full_adder fa91(.a(weight_0_12[9]), .b(weight_0_12[10]), .cin(weight_0_12[11]), .sum(weight_1_12[7]), .cout(weight_1_13[6]));
full_adder fa92(.a(weight_0_13[9]), .b(weight_0_13[10]), .cin(weight_0_13[11]), .sum(weight_1_13[7]), .cout(weight_1_14[6]));
full_adder fa93(.a(weight_0_14[9]), .b(weight_0_14[10]), .cin(weight_0_14[11]), .sum(weight_1_14[7]), .cout(weight_1_15[6]));
full_adder fa94(.a(weight_0_15[9]), .b(weight_0_15[10]), .cin(weight_0_15[11]), .sum(weight_1_15[7]), .cout(weight_1_16[6]));
full_adder fa95(.a(weight_0_16[9]), .b(weight_0_16[10]), .cin(weight_0_16[11]), .sum(weight_1_16[7]), .cout(weight_1_17[6]));
full_adder fa96(.a(weight_0_17[9]), .b(weight_0_17[10]), .cin(weight_0_17[11]), .sum(weight_1_17[7]), .cout(weight_1_18[6]));
full_adder fa97(.a(weight_0_18[9]), .b(weight_0_18[10]), .cin(weight_0_18[11]), .sum(weight_1_18[7]), .cout(weight_1_19[6]));
full_adder fa98(.a(weight_0_19[9]), .b(weight_0_19[10]), .cin(weight_0_19[11]), .sum(weight_1_19[7]), .cout(weight_1_20[6]));
full_adder fa99(.a(weight_0_20[9]), .b(weight_0_20[10]), .cin(weight_0_20[11]), .sum(weight_1_20[7]), .cout(weight_1_21[6]));
full_adder fa100(.a(weight_0_21[9]), .b(weight_0_21[10]), .cin(weight_0_21[11]), .sum(weight_1_21[7]), .cout(weight_1_22[6]));
full_adder fa101(.a(weight_0_22[9]), .b(weight_0_22[10]), .cin(weight_0_22[11]), .sum(weight_1_22[7]), .cout(weight_1_23[6]));
full_adder fa102(.a(weight_0_23[9]), .b(weight_0_23[10]), .cin(weight_0_23[11]), .sum(weight_1_23[7]), .cout(weight_1_24[6]));
full_adder fa103(.a(weight_0_24[9]), .b(weight_0_24[10]), .cin(weight_0_24[11]), .sum(weight_1_24[7]), .cout(weight_1_25[6]));
full_adder fa104(.a(weight_0_25[9]), .b(weight_0_25[10]), .cin(weight_0_25[11]), .sum(weight_1_25[7]), .cout(weight_1_26[6]));
full_adder fa105(.a(weight_0_26[9]), .b(weight_0_26[10]), .cin(weight_0_26[11]), .sum(weight_1_26[7]), .cout(weight_1_27[6]));
full_adder fa106(.a(weight_0_27[9]), .b(weight_0_27[10]), .cin(weight_0_27[11]), .sum(weight_1_27[7]), .cout(weight_1_28[6]));
full_adder fa107(.a(weight_0_28[9]), .b(weight_0_28[10]), .cin(weight_0_28[11]), .sum(weight_1_28[7]), .cout(weight_1_29[6]));
full_adder fa108(.a(weight_0_29[9]), .b(weight_0_29[10]), .cin(weight_0_29[11]), .sum(weight_1_29[7]), .cout(weight_1_30[6]));
full_adder fa109(.a(weight_0_30[9]), .b(weight_0_30[10]), .cin(weight_0_30[11]), .sum(weight_1_30[7]), .cout(weight_1_31[6]));
full_adder fa110(.a(weight_0_31[9]), .b(weight_0_31[10]), .cin(weight_0_31[11]), .sum(weight_1_31[7]), .cout(weight_1_32[6]));
full_adder fa111(.a(weight_0_32[8]), .b(weight_0_32[9]), .cin(weight_0_32[10]), .sum(weight_1_32[7]), .cout(weight_1_33[6]));
full_adder fa112(.a(weight_0_33[7]), .b(weight_0_33[8]), .cin(weight_0_33[9]), .sum(weight_1_33[7]), .cout(weight_1_34[4]));
full_adder fa113(.a(weight_0_34[6]), .b(weight_0_34[7]), .cin(weight_0_34[8]), .sum(weight_1_34[5]), .cout(weight_1_35[4]));
full_adder fa114(.a(weight_0_35[5]), .b(weight_0_35[6]), .cin(weight_0_35[7]), .sum(weight_1_35[5]), .cout(weight_1_36[4]));
full_adder fa115(.a(weight_0_36[4]), .b(weight_0_36[5]), .cin(weight_0_36[6]), .sum(weight_1_36[5]), .cout(weight_1_37[2]));
full_adder fa116(.a(weight_0_37[3]), .b(weight_0_37[4]), .cin(weight_0_37[5]), .sum(weight_1_37[3]), .cout(weight_1_38[2]));
full_adder fa117(.a(weight_0_38[2]), .b(weight_0_38[3]), .cin(weight_0_38[4]), .sum(weight_1_38[3]), .cout(weight_1_39[2]));
full_adder fa118(.a(weight_0_39[1]), .b(weight_0_39[2]), .cin(weight_0_39[3]), .sum(weight_1_39[3]), .cout(weight_1_40[0]));
full_adder fa119(.a(weight_0_40[0]), .b(weight_0_40[1]), .cin(weight_0_40[2]), .sum(weight_1_40[1]), .cout(weight_1_41[0]));
half_adder ha7(.a(weight_0_41[0]), .b(weight_0_41[1]), .sum(weight_1_41[1]), .cout(weight_1_42[0]));
assign weight_1_42[1] = weight_0_42[0];
assign weight_1_12[8] = weight_0_12[12];
half_adder ha8(.a(weight_0_13[12]), .b(weight_0_13[13]), .sum(weight_1_13[8]), .cout(weight_1_14[8]));
full_adder fa120(.a(weight_0_14[12]), .b(weight_0_14[13]), .cin(weight_0_14[14]), .sum(weight_1_14[9]), .cout(weight_1_15[8]));
full_adder fa121(.a(weight_0_15[12]), .b(weight_0_15[13]), .cin(weight_0_15[14]), .sum(weight_1_15[9]), .cout(weight_1_16[8]));
full_adder fa122(.a(weight_0_16[12]), .b(weight_0_16[13]), .cin(weight_0_16[14]), .sum(weight_1_16[9]), .cout(weight_1_17[8]));
full_adder fa123(.a(weight_0_17[12]), .b(weight_0_17[13]), .cin(weight_0_17[14]), .sum(weight_1_17[9]), .cout(weight_1_18[8]));
full_adder fa124(.a(weight_0_18[12]), .b(weight_0_18[13]), .cin(weight_0_18[14]), .sum(weight_1_18[9]), .cout(weight_1_19[8]));
full_adder fa125(.a(weight_0_19[12]), .b(weight_0_19[13]), .cin(weight_0_19[14]), .sum(weight_1_19[9]), .cout(weight_1_20[8]));
full_adder fa126(.a(weight_0_20[12]), .b(weight_0_20[13]), .cin(weight_0_20[14]), .sum(weight_1_20[9]), .cout(weight_1_21[8]));
full_adder fa127(.a(weight_0_21[12]), .b(weight_0_21[13]), .cin(weight_0_21[14]), .sum(weight_1_21[9]), .cout(weight_1_22[8]));
full_adder fa128(.a(weight_0_22[12]), .b(weight_0_22[13]), .cin(weight_0_22[14]), .sum(weight_1_22[9]), .cout(weight_1_23[8]));
full_adder fa129(.a(weight_0_23[12]), .b(weight_0_23[13]), .cin(weight_0_23[14]), .sum(weight_1_23[9]), .cout(weight_1_24[8]));
full_adder fa130(.a(weight_0_24[12]), .b(weight_0_24[13]), .cin(weight_0_24[14]), .sum(weight_1_24[9]), .cout(weight_1_25[8]));
full_adder fa131(.a(weight_0_25[12]), .b(weight_0_25[13]), .cin(weight_0_25[14]), .sum(weight_1_25[9]), .cout(weight_1_26[8]));
full_adder fa132(.a(weight_0_26[12]), .b(weight_0_26[13]), .cin(weight_0_26[14]), .sum(weight_1_26[9]), .cout(weight_1_27[8]));
full_adder fa133(.a(weight_0_27[12]), .b(weight_0_27[13]), .cin(weight_0_27[14]), .sum(weight_1_27[9]), .cout(weight_1_28[8]));
full_adder fa134(.a(weight_0_28[12]), .b(weight_0_28[13]), .cin(weight_0_28[14]), .sum(weight_1_28[9]), .cout(weight_1_29[8]));
full_adder fa135(.a(weight_0_29[12]), .b(weight_0_29[13]), .cin(weight_0_29[14]), .sum(weight_1_29[9]), .cout(weight_1_30[8]));
full_adder fa136(.a(weight_0_30[12]), .b(weight_0_30[13]), .cin(weight_0_30[14]), .sum(weight_1_30[9]), .cout(weight_1_31[8]));
full_adder fa137(.a(weight_0_31[12]), .b(weight_0_31[13]), .cin(weight_0_31[14]), .sum(weight_1_31[9]), .cout(weight_1_32[8]));
full_adder fa138(.a(weight_0_32[11]), .b(weight_0_32[12]), .cin(weight_0_32[13]), .sum(weight_1_32[9]), .cout(weight_1_33[8]));
full_adder fa139(.a(weight_0_33[10]), .b(weight_0_33[11]), .cin(weight_0_33[12]), .sum(weight_1_33[9]), .cout(weight_1_34[6]));
full_adder fa140(.a(weight_0_34[9]), .b(weight_0_34[10]), .cin(weight_0_34[11]), .sum(weight_1_34[7]), .cout(weight_1_35[6]));
full_adder fa141(.a(weight_0_35[8]), .b(weight_0_35[9]), .cin(weight_0_35[10]), .sum(weight_1_35[7]), .cout(weight_1_36[6]));
full_adder fa142(.a(weight_0_36[7]), .b(weight_0_36[8]), .cin(weight_0_36[9]), .sum(weight_1_36[7]), .cout(weight_1_37[4]));
full_adder fa143(.a(weight_0_37[6]), .b(weight_0_37[7]), .cin(weight_0_37[8]), .sum(weight_1_37[5]), .cout(weight_1_38[4]));
full_adder fa144(.a(weight_0_38[5]), .b(weight_0_38[6]), .cin(weight_0_38[7]), .sum(weight_1_38[5]), .cout(weight_1_39[4]));
full_adder fa145(.a(weight_0_39[4]), .b(weight_0_39[5]), .cin(weight_0_39[6]), .sum(weight_1_39[5]), .cout(weight_1_40[2]));
full_adder fa146(.a(weight_0_40[3]), .b(weight_0_40[4]), .cin(weight_0_40[5]), .sum(weight_1_40[3]), .cout(weight_1_41[2]));
full_adder fa147(.a(weight_0_41[2]), .b(weight_0_41[3]), .cin(weight_0_41[4]), .sum(weight_1_41[3]), .cout(weight_1_42[2]));
full_adder fa148(.a(weight_0_42[1]), .b(weight_0_42[2]), .cin(weight_0_42[3]), .sum(weight_1_42[3]), .cout(weight_1_43[0]));
full_adder fa149(.a(weight_0_43[0]), .b(weight_0_43[1]), .cin(weight_0_43[2]), .sum(weight_1_43[1]), .cout(weight_1_44[0]));
half_adder ha9(.a(weight_0_44[0]), .b(weight_0_44[1]), .sum(weight_1_44[1]), .cout(weight_1_45[0]));
assign weight_1_45[1] = weight_0_45[0];
assign weight_1_15[10] = weight_0_15[15];
half_adder ha10(.a(weight_0_16[15]), .b(weight_0_16[16]), .sum(weight_1_16[10]), .cout(weight_1_17[10]));
full_adder fa150(.a(weight_0_17[15]), .b(weight_0_17[16]), .cin(weight_0_17[17]), .sum(weight_1_17[11]), .cout(weight_1_18[10]));
full_adder fa151(.a(weight_0_18[15]), .b(weight_0_18[16]), .cin(weight_0_18[17]), .sum(weight_1_18[11]), .cout(weight_1_19[10]));
full_adder fa152(.a(weight_0_19[15]), .b(weight_0_19[16]), .cin(weight_0_19[17]), .sum(weight_1_19[11]), .cout(weight_1_20[10]));
full_adder fa153(.a(weight_0_20[15]), .b(weight_0_20[16]), .cin(weight_0_20[17]), .sum(weight_1_20[11]), .cout(weight_1_21[10]));
full_adder fa154(.a(weight_0_21[15]), .b(weight_0_21[16]), .cin(weight_0_21[17]), .sum(weight_1_21[11]), .cout(weight_1_22[10]));
full_adder fa155(.a(weight_0_22[15]), .b(weight_0_22[16]), .cin(weight_0_22[17]), .sum(weight_1_22[11]), .cout(weight_1_23[10]));
full_adder fa156(.a(weight_0_23[15]), .b(weight_0_23[16]), .cin(weight_0_23[17]), .sum(weight_1_23[11]), .cout(weight_1_24[10]));
full_adder fa157(.a(weight_0_24[15]), .b(weight_0_24[16]), .cin(weight_0_24[17]), .sum(weight_1_24[11]), .cout(weight_1_25[10]));
full_adder fa158(.a(weight_0_25[15]), .b(weight_0_25[16]), .cin(weight_0_25[17]), .sum(weight_1_25[11]), .cout(weight_1_26[10]));
full_adder fa159(.a(weight_0_26[15]), .b(weight_0_26[16]), .cin(weight_0_26[17]), .sum(weight_1_26[11]), .cout(weight_1_27[10]));
full_adder fa160(.a(weight_0_27[15]), .b(weight_0_27[16]), .cin(weight_0_27[17]), .sum(weight_1_27[11]), .cout(weight_1_28[10]));
full_adder fa161(.a(weight_0_28[15]), .b(weight_0_28[16]), .cin(weight_0_28[17]), .sum(weight_1_28[11]), .cout(weight_1_29[10]));
full_adder fa162(.a(weight_0_29[15]), .b(weight_0_29[16]), .cin(weight_0_29[17]), .sum(weight_1_29[11]), .cout(weight_1_30[10]));
full_adder fa163(.a(weight_0_30[15]), .b(weight_0_30[16]), .cin(weight_0_30[17]), .sum(weight_1_30[11]), .cout(weight_1_31[10]));
full_adder fa164(.a(weight_0_31[15]), .b(weight_0_31[16]), .cin(weight_0_31[17]), .sum(weight_1_31[11]), .cout(weight_1_32[10]));
full_adder fa165(.a(weight_0_32[14]), .b(weight_0_32[15]), .cin(weight_0_32[16]), .sum(weight_1_32[11]), .cout(weight_1_33[10]));
full_adder fa166(.a(weight_0_33[13]), .b(weight_0_33[14]), .cin(weight_0_33[15]), .sum(weight_1_33[11]), .cout(weight_1_34[8]));
full_adder fa167(.a(weight_0_34[12]), .b(weight_0_34[13]), .cin(weight_0_34[14]), .sum(weight_1_34[9]), .cout(weight_1_35[8]));
full_adder fa168(.a(weight_0_35[11]), .b(weight_0_35[12]), .cin(weight_0_35[13]), .sum(weight_1_35[9]), .cout(weight_1_36[8]));
full_adder fa169(.a(weight_0_36[10]), .b(weight_0_36[11]), .cin(weight_0_36[12]), .sum(weight_1_36[9]), .cout(weight_1_37[6]));
full_adder fa170(.a(weight_0_37[9]), .b(weight_0_37[10]), .cin(weight_0_37[11]), .sum(weight_1_37[7]), .cout(weight_1_38[6]));
full_adder fa171(.a(weight_0_38[8]), .b(weight_0_38[9]), .cin(weight_0_38[10]), .sum(weight_1_38[7]), .cout(weight_1_39[6]));
full_adder fa172(.a(weight_0_39[7]), .b(weight_0_39[8]), .cin(weight_0_39[9]), .sum(weight_1_39[7]), .cout(weight_1_40[4]));
full_adder fa173(.a(weight_0_40[6]), .b(weight_0_40[7]), .cin(weight_0_40[8]), .sum(weight_1_40[5]), .cout(weight_1_41[4]));
full_adder fa174(.a(weight_0_41[5]), .b(weight_0_41[6]), .cin(weight_0_41[7]), .sum(weight_1_41[5]), .cout(weight_1_42[4]));
full_adder fa175(.a(weight_0_42[4]), .b(weight_0_42[5]), .cin(weight_0_42[6]), .sum(weight_1_42[5]), .cout(weight_1_43[2]));
full_adder fa176(.a(weight_0_43[3]), .b(weight_0_43[4]), .cin(weight_0_43[5]), .sum(weight_1_43[3]), .cout(weight_1_44[2]));
full_adder fa177(.a(weight_0_44[2]), .b(weight_0_44[3]), .cin(weight_0_44[4]), .sum(weight_1_44[3]), .cout(weight_1_45[2]));
full_adder fa178(.a(weight_0_45[1]), .b(weight_0_45[2]), .cin(weight_0_45[3]), .sum(weight_1_45[3]), .cout(weight_1_46[0]));
full_adder fa179(.a(weight_0_46[0]), .b(weight_0_46[1]), .cin(weight_0_46[2]), .sum(weight_1_46[1]), .cout(weight_1_47[0]));
half_adder ha11(.a(weight_0_47[0]), .b(weight_0_47[1]), .sum(weight_1_47[1]), .cout(weight_1_48[0]));
assign weight_1_48[1] = weight_0_48[0];
assign weight_1_18[12] = weight_0_18[18];
half_adder ha12(.a(weight_0_19[18]), .b(weight_0_19[19]), .sum(weight_1_19[12]), .cout(weight_1_20[12]));
full_adder fa180(.a(weight_0_20[18]), .b(weight_0_20[19]), .cin(weight_0_20[20]), .sum(weight_1_20[13]), .cout(weight_1_21[12]));
full_adder fa181(.a(weight_0_21[18]), .b(weight_0_21[19]), .cin(weight_0_21[20]), .sum(weight_1_21[13]), .cout(weight_1_22[12]));
full_adder fa182(.a(weight_0_22[18]), .b(weight_0_22[19]), .cin(weight_0_22[20]), .sum(weight_1_22[13]), .cout(weight_1_23[12]));
full_adder fa183(.a(weight_0_23[18]), .b(weight_0_23[19]), .cin(weight_0_23[20]), .sum(weight_1_23[13]), .cout(weight_1_24[12]));
full_adder fa184(.a(weight_0_24[18]), .b(weight_0_24[19]), .cin(weight_0_24[20]), .sum(weight_1_24[13]), .cout(weight_1_25[12]));
full_adder fa185(.a(weight_0_25[18]), .b(weight_0_25[19]), .cin(weight_0_25[20]), .sum(weight_1_25[13]), .cout(weight_1_26[12]));
full_adder fa186(.a(weight_0_26[18]), .b(weight_0_26[19]), .cin(weight_0_26[20]), .sum(weight_1_26[13]), .cout(weight_1_27[12]));
full_adder fa187(.a(weight_0_27[18]), .b(weight_0_27[19]), .cin(weight_0_27[20]), .sum(weight_1_27[13]), .cout(weight_1_28[12]));
full_adder fa188(.a(weight_0_28[18]), .b(weight_0_28[19]), .cin(weight_0_28[20]), .sum(weight_1_28[13]), .cout(weight_1_29[12]));
full_adder fa189(.a(weight_0_29[18]), .b(weight_0_29[19]), .cin(weight_0_29[20]), .sum(weight_1_29[13]), .cout(weight_1_30[12]));
full_adder fa190(.a(weight_0_30[18]), .b(weight_0_30[19]), .cin(weight_0_30[20]), .sum(weight_1_30[13]), .cout(weight_1_31[12]));
full_adder fa191(.a(weight_0_31[18]), .b(weight_0_31[19]), .cin(weight_0_31[20]), .sum(weight_1_31[13]), .cout(weight_1_32[12]));
full_adder fa192(.a(weight_0_32[17]), .b(weight_0_32[18]), .cin(weight_0_32[19]), .sum(weight_1_32[13]), .cout(weight_1_33[12]));
full_adder fa193(.a(weight_0_33[16]), .b(weight_0_33[17]), .cin(weight_0_33[18]), .sum(weight_1_33[13]), .cout(weight_1_34[10]));
full_adder fa194(.a(weight_0_34[15]), .b(weight_0_34[16]), .cin(weight_0_34[17]), .sum(weight_1_34[11]), .cout(weight_1_35[10]));
full_adder fa195(.a(weight_0_35[14]), .b(weight_0_35[15]), .cin(weight_0_35[16]), .sum(weight_1_35[11]), .cout(weight_1_36[10]));
full_adder fa196(.a(weight_0_36[13]), .b(weight_0_36[14]), .cin(weight_0_36[15]), .sum(weight_1_36[11]), .cout(weight_1_37[8]));
full_adder fa197(.a(weight_0_37[12]), .b(weight_0_37[13]), .cin(weight_0_37[14]), .sum(weight_1_37[9]), .cout(weight_1_38[8]));
full_adder fa198(.a(weight_0_38[11]), .b(weight_0_38[12]), .cin(weight_0_38[13]), .sum(weight_1_38[9]), .cout(weight_1_39[8]));
full_adder fa199(.a(weight_0_39[10]), .b(weight_0_39[11]), .cin(weight_0_39[12]), .sum(weight_1_39[9]), .cout(weight_1_40[6]));
full_adder fa200(.a(weight_0_40[9]), .b(weight_0_40[10]), .cin(weight_0_40[11]), .sum(weight_1_40[7]), .cout(weight_1_41[6]));
full_adder fa201(.a(weight_0_41[8]), .b(weight_0_41[9]), .cin(weight_0_41[10]), .sum(weight_1_41[7]), .cout(weight_1_42[6]));
full_adder fa202(.a(weight_0_42[7]), .b(weight_0_42[8]), .cin(weight_0_42[9]), .sum(weight_1_42[7]), .cout(weight_1_43[4]));
full_adder fa203(.a(weight_0_43[6]), .b(weight_0_43[7]), .cin(weight_0_43[8]), .sum(weight_1_43[5]), .cout(weight_1_44[4]));
full_adder fa204(.a(weight_0_44[5]), .b(weight_0_44[6]), .cin(weight_0_44[7]), .sum(weight_1_44[5]), .cout(weight_1_45[4]));
full_adder fa205(.a(weight_0_45[4]), .b(weight_0_45[5]), .cin(weight_0_45[6]), .sum(weight_1_45[5]), .cout(weight_1_46[2]));
full_adder fa206(.a(weight_0_46[3]), .b(weight_0_46[4]), .cin(weight_0_46[5]), .sum(weight_1_46[3]), .cout(weight_1_47[2]));
full_adder fa207(.a(weight_0_47[2]), .b(weight_0_47[3]), .cin(weight_0_47[4]), .sum(weight_1_47[3]), .cout(weight_1_48[2]));
full_adder fa208(.a(weight_0_48[1]), .b(weight_0_48[2]), .cin(weight_0_48[3]), .sum(weight_1_48[3]), .cout(weight_1_49[0]));
full_adder fa209(.a(weight_0_49[0]), .b(weight_0_49[1]), .cin(weight_0_49[2]), .sum(weight_1_49[1]), .cout(weight_1_50[0]));
half_adder ha13(.a(weight_0_50[0]), .b(weight_0_50[1]), .sum(weight_1_50[1]), .cout(weight_1_51[0]));
assign weight_1_51[1] = weight_0_51[0];
assign weight_1_21[14] = weight_0_21[21];
half_adder ha14(.a(weight_0_22[21]), .b(weight_0_22[22]), .sum(weight_1_22[14]), .cout(weight_1_23[14]));
full_adder fa210(.a(weight_0_23[21]), .b(weight_0_23[22]), .cin(weight_0_23[23]), .sum(weight_1_23[15]), .cout(weight_1_24[14]));
full_adder fa211(.a(weight_0_24[21]), .b(weight_0_24[22]), .cin(weight_0_24[23]), .sum(weight_1_24[15]), .cout(weight_1_25[14]));
full_adder fa212(.a(weight_0_25[21]), .b(weight_0_25[22]), .cin(weight_0_25[23]), .sum(weight_1_25[15]), .cout(weight_1_26[14]));
full_adder fa213(.a(weight_0_26[21]), .b(weight_0_26[22]), .cin(weight_0_26[23]), .sum(weight_1_26[15]), .cout(weight_1_27[14]));
full_adder fa214(.a(weight_0_27[21]), .b(weight_0_27[22]), .cin(weight_0_27[23]), .sum(weight_1_27[15]), .cout(weight_1_28[14]));
full_adder fa215(.a(weight_0_28[21]), .b(weight_0_28[22]), .cin(weight_0_28[23]), .sum(weight_1_28[15]), .cout(weight_1_29[14]));
full_adder fa216(.a(weight_0_29[21]), .b(weight_0_29[22]), .cin(weight_0_29[23]), .sum(weight_1_29[15]), .cout(weight_1_30[14]));
full_adder fa217(.a(weight_0_30[21]), .b(weight_0_30[22]), .cin(weight_0_30[23]), .sum(weight_1_30[15]), .cout(weight_1_31[14]));
full_adder fa218(.a(weight_0_31[21]), .b(weight_0_31[22]), .cin(weight_0_31[23]), .sum(weight_1_31[15]), .cout(weight_1_32[14]));
full_adder fa219(.a(weight_0_32[20]), .b(weight_0_32[21]), .cin(weight_0_32[22]), .sum(weight_1_32[15]), .cout(weight_1_33[14]));
full_adder fa220(.a(weight_0_33[19]), .b(weight_0_33[20]), .cin(weight_0_33[21]), .sum(weight_1_33[15]), .cout(weight_1_34[12]));
full_adder fa221(.a(weight_0_34[18]), .b(weight_0_34[19]), .cin(weight_0_34[20]), .sum(weight_1_34[13]), .cout(weight_1_35[12]));
full_adder fa222(.a(weight_0_35[17]), .b(weight_0_35[18]), .cin(weight_0_35[19]), .sum(weight_1_35[13]), .cout(weight_1_36[12]));
full_adder fa223(.a(weight_0_36[16]), .b(weight_0_36[17]), .cin(weight_0_36[18]), .sum(weight_1_36[13]), .cout(weight_1_37[10]));
full_adder fa224(.a(weight_0_37[15]), .b(weight_0_37[16]), .cin(weight_0_37[17]), .sum(weight_1_37[11]), .cout(weight_1_38[10]));
full_adder fa225(.a(weight_0_38[14]), .b(weight_0_38[15]), .cin(weight_0_38[16]), .sum(weight_1_38[11]), .cout(weight_1_39[10]));
full_adder fa226(.a(weight_0_39[13]), .b(weight_0_39[14]), .cin(weight_0_39[15]), .sum(weight_1_39[11]), .cout(weight_1_40[8]));
full_adder fa227(.a(weight_0_40[12]), .b(weight_0_40[13]), .cin(weight_0_40[14]), .sum(weight_1_40[9]), .cout(weight_1_41[8]));
full_adder fa228(.a(weight_0_41[11]), .b(weight_0_41[12]), .cin(weight_0_41[13]), .sum(weight_1_41[9]), .cout(weight_1_42[8]));
full_adder fa229(.a(weight_0_42[10]), .b(weight_0_42[11]), .cin(weight_0_42[12]), .sum(weight_1_42[9]), .cout(weight_1_43[6]));
full_adder fa230(.a(weight_0_43[9]), .b(weight_0_43[10]), .cin(weight_0_43[11]), .sum(weight_1_43[7]), .cout(weight_1_44[6]));
full_adder fa231(.a(weight_0_44[8]), .b(weight_0_44[9]), .cin(weight_0_44[10]), .sum(weight_1_44[7]), .cout(weight_1_45[6]));
full_adder fa232(.a(weight_0_45[7]), .b(weight_0_45[8]), .cin(weight_0_45[9]), .sum(weight_1_45[7]), .cout(weight_1_46[4]));
full_adder fa233(.a(weight_0_46[6]), .b(weight_0_46[7]), .cin(weight_0_46[8]), .sum(weight_1_46[5]), .cout(weight_1_47[4]));
full_adder fa234(.a(weight_0_47[5]), .b(weight_0_47[6]), .cin(weight_0_47[7]), .sum(weight_1_47[5]), .cout(weight_1_48[4]));
full_adder fa235(.a(weight_0_48[4]), .b(weight_0_48[5]), .cin(weight_0_48[6]), .sum(weight_1_48[5]), .cout(weight_1_49[2]));
full_adder fa236(.a(weight_0_49[3]), .b(weight_0_49[4]), .cin(weight_0_49[5]), .sum(weight_1_49[3]), .cout(weight_1_50[2]));
full_adder fa237(.a(weight_0_50[2]), .b(weight_0_50[3]), .cin(weight_0_50[4]), .sum(weight_1_50[3]), .cout(weight_1_51[2]));
full_adder fa238(.a(weight_0_51[1]), .b(weight_0_51[2]), .cin(weight_0_51[3]), .sum(weight_1_51[3]), .cout(weight_1_52[0]));
full_adder fa239(.a(weight_0_52[0]), .b(weight_0_52[1]), .cin(weight_0_52[2]), .sum(weight_1_52[1]), .cout(weight_1_53[0]));
half_adder ha15(.a(weight_0_53[0]), .b(weight_0_53[1]), .sum(weight_1_53[1]), .cout(weight_1_54[0]));
assign weight_1_54[1] = weight_0_54[0];
assign weight_1_24[16] = weight_0_24[24];
half_adder ha16(.a(weight_0_25[24]), .b(weight_0_25[25]), .sum(weight_1_25[16]), .cout(weight_1_26[16]));
full_adder fa240(.a(weight_0_26[24]), .b(weight_0_26[25]), .cin(weight_0_26[26]), .sum(weight_1_26[17]), .cout(weight_1_27[16]));
full_adder fa241(.a(weight_0_27[24]), .b(weight_0_27[25]), .cin(weight_0_27[26]), .sum(weight_1_27[17]), .cout(weight_1_28[16]));
full_adder fa242(.a(weight_0_28[24]), .b(weight_0_28[25]), .cin(weight_0_28[26]), .sum(weight_1_28[17]), .cout(weight_1_29[16]));
full_adder fa243(.a(weight_0_29[24]), .b(weight_0_29[25]), .cin(weight_0_29[26]), .sum(weight_1_29[17]), .cout(weight_1_30[16]));
full_adder fa244(.a(weight_0_30[24]), .b(weight_0_30[25]), .cin(weight_0_30[26]), .sum(weight_1_30[17]), .cout(weight_1_31[16]));
full_adder fa245(.a(weight_0_31[24]), .b(weight_0_31[25]), .cin(weight_0_31[26]), .sum(weight_1_31[17]), .cout(weight_1_32[16]));
full_adder fa246(.a(weight_0_32[23]), .b(weight_0_32[24]), .cin(weight_0_32[25]), .sum(weight_1_32[17]), .cout(weight_1_33[16]));
full_adder fa247(.a(weight_0_33[22]), .b(weight_0_33[23]), .cin(weight_0_33[24]), .sum(weight_1_33[17]), .cout(weight_1_34[14]));
full_adder fa248(.a(weight_0_34[21]), .b(weight_0_34[22]), .cin(weight_0_34[23]), .sum(weight_1_34[15]), .cout(weight_1_35[14]));
full_adder fa249(.a(weight_0_35[20]), .b(weight_0_35[21]), .cin(weight_0_35[22]), .sum(weight_1_35[15]), .cout(weight_1_36[14]));
full_adder fa250(.a(weight_0_36[19]), .b(weight_0_36[20]), .cin(weight_0_36[21]), .sum(weight_1_36[15]), .cout(weight_1_37[12]));
full_adder fa251(.a(weight_0_37[18]), .b(weight_0_37[19]), .cin(weight_0_37[20]), .sum(weight_1_37[13]), .cout(weight_1_38[12]));
full_adder fa252(.a(weight_0_38[17]), .b(weight_0_38[18]), .cin(weight_0_38[19]), .sum(weight_1_38[13]), .cout(weight_1_39[12]));
full_adder fa253(.a(weight_0_39[16]), .b(weight_0_39[17]), .cin(weight_0_39[18]), .sum(weight_1_39[13]), .cout(weight_1_40[10]));
full_adder fa254(.a(weight_0_40[15]), .b(weight_0_40[16]), .cin(weight_0_40[17]), .sum(weight_1_40[11]), .cout(weight_1_41[10]));
full_adder fa255(.a(weight_0_41[14]), .b(weight_0_41[15]), .cin(weight_0_41[16]), .sum(weight_1_41[11]), .cout(weight_1_42[10]));
full_adder fa256(.a(weight_0_42[13]), .b(weight_0_42[14]), .cin(weight_0_42[15]), .sum(weight_1_42[11]), .cout(weight_1_43[8]));
full_adder fa257(.a(weight_0_43[12]), .b(weight_0_43[13]), .cin(weight_0_43[14]), .sum(weight_1_43[9]), .cout(weight_1_44[8]));
full_adder fa258(.a(weight_0_44[11]), .b(weight_0_44[12]), .cin(weight_0_44[13]), .sum(weight_1_44[9]), .cout(weight_1_45[8]));
full_adder fa259(.a(weight_0_45[10]), .b(weight_0_45[11]), .cin(weight_0_45[12]), .sum(weight_1_45[9]), .cout(weight_1_46[6]));
full_adder fa260(.a(weight_0_46[9]), .b(weight_0_46[10]), .cin(weight_0_46[11]), .sum(weight_1_46[7]), .cout(weight_1_47[6]));
full_adder fa261(.a(weight_0_47[8]), .b(weight_0_47[9]), .cin(weight_0_47[10]), .sum(weight_1_47[7]), .cout(weight_1_48[6]));
full_adder fa262(.a(weight_0_48[7]), .b(weight_0_48[8]), .cin(weight_0_48[9]), .sum(weight_1_48[7]), .cout(weight_1_49[4]));
full_adder fa263(.a(weight_0_49[6]), .b(weight_0_49[7]), .cin(weight_0_49[8]), .sum(weight_1_49[5]), .cout(weight_1_50[4]));
full_adder fa264(.a(weight_0_50[5]), .b(weight_0_50[6]), .cin(weight_0_50[7]), .sum(weight_1_50[5]), .cout(weight_1_51[4]));
full_adder fa265(.a(weight_0_51[4]), .b(weight_0_51[5]), .cin(weight_0_51[6]), .sum(weight_1_51[5]), .cout(weight_1_52[2]));
full_adder fa266(.a(weight_0_52[3]), .b(weight_0_52[4]), .cin(weight_0_52[5]), .sum(weight_1_52[3]), .cout(weight_1_53[2]));
full_adder fa267(.a(weight_0_53[2]), .b(weight_0_53[3]), .cin(weight_0_53[4]), .sum(weight_1_53[3]), .cout(weight_1_54[2]));
full_adder fa268(.a(weight_0_54[1]), .b(weight_0_54[2]), .cin(weight_0_54[3]), .sum(weight_1_54[3]), .cout(weight_1_55[0]));
full_adder fa269(.a(weight_0_55[0]), .b(weight_0_55[1]), .cin(weight_0_55[2]), .sum(weight_1_55[1]), .cout(weight_1_56[0]));
half_adder ha17(.a(weight_0_56[0]), .b(weight_0_56[1]), .sum(weight_1_56[1]), .cout(weight_1_57[0]));
assign weight_1_57[1] = weight_0_57[0];
assign weight_1_27[18] = weight_0_27[27];
half_adder ha18(.a(weight_0_28[27]), .b(weight_0_28[28]), .sum(weight_1_28[18]), .cout(weight_1_29[18]));
full_adder fa270(.a(weight_0_29[27]), .b(weight_0_29[28]), .cin(weight_0_29[29]), .sum(weight_1_29[19]), .cout(weight_1_30[18]));
full_adder fa271(.a(weight_0_30[27]), .b(weight_0_30[28]), .cin(weight_0_30[29]), .sum(weight_1_30[19]), .cout(weight_1_31[18]));
full_adder fa272(.a(weight_0_31[27]), .b(weight_0_31[28]), .cin(weight_0_31[29]), .sum(weight_1_31[19]), .cout(weight_1_32[18]));
full_adder fa273(.a(weight_0_32[26]), .b(weight_0_32[27]), .cin(weight_0_32[28]), .sum(weight_1_32[19]), .cout(weight_1_33[18]));
full_adder fa274(.a(weight_0_33[25]), .b(weight_0_33[26]), .cin(weight_0_33[27]), .sum(weight_1_33[19]), .cout(weight_1_34[16]));
full_adder fa275(.a(weight_0_34[24]), .b(weight_0_34[25]), .cin(weight_0_34[26]), .sum(weight_1_34[17]), .cout(weight_1_35[16]));
full_adder fa276(.a(weight_0_35[23]), .b(weight_0_35[24]), .cin(weight_0_35[25]), .sum(weight_1_35[17]), .cout(weight_1_36[16]));
full_adder fa277(.a(weight_0_36[22]), .b(weight_0_36[23]), .cin(weight_0_36[24]), .sum(weight_1_36[17]), .cout(weight_1_37[14]));
full_adder fa278(.a(weight_0_37[21]), .b(weight_0_37[22]), .cin(weight_0_37[23]), .sum(weight_1_37[15]), .cout(weight_1_38[14]));
full_adder fa279(.a(weight_0_38[20]), .b(weight_0_38[21]), .cin(weight_0_38[22]), .sum(weight_1_38[15]), .cout(weight_1_39[14]));
full_adder fa280(.a(weight_0_39[19]), .b(weight_0_39[20]), .cin(weight_0_39[21]), .sum(weight_1_39[15]), .cout(weight_1_40[12]));
full_adder fa281(.a(weight_0_40[18]), .b(weight_0_40[19]), .cin(weight_0_40[20]), .sum(weight_1_40[13]), .cout(weight_1_41[12]));
full_adder fa282(.a(weight_0_41[17]), .b(weight_0_41[18]), .cin(weight_0_41[19]), .sum(weight_1_41[13]), .cout(weight_1_42[12]));
full_adder fa283(.a(weight_0_42[16]), .b(weight_0_42[17]), .cin(weight_0_42[18]), .sum(weight_1_42[13]), .cout(weight_1_43[10]));
full_adder fa284(.a(weight_0_43[15]), .b(weight_0_43[16]), .cin(weight_0_43[17]), .sum(weight_1_43[11]), .cout(weight_1_44[10]));
full_adder fa285(.a(weight_0_44[14]), .b(weight_0_44[15]), .cin(weight_0_44[16]), .sum(weight_1_44[11]), .cout(weight_1_45[10]));
full_adder fa286(.a(weight_0_45[13]), .b(weight_0_45[14]), .cin(weight_0_45[15]), .sum(weight_1_45[11]), .cout(weight_1_46[8]));
full_adder fa287(.a(weight_0_46[12]), .b(weight_0_46[13]), .cin(weight_0_46[14]), .sum(weight_1_46[9]), .cout(weight_1_47[8]));
full_adder fa288(.a(weight_0_47[11]), .b(weight_0_47[12]), .cin(weight_0_47[13]), .sum(weight_1_47[9]), .cout(weight_1_48[8]));
full_adder fa289(.a(weight_0_48[10]), .b(weight_0_48[11]), .cin(weight_0_48[12]), .sum(weight_1_48[9]), .cout(weight_1_49[6]));
full_adder fa290(.a(weight_0_49[9]), .b(weight_0_49[10]), .cin(weight_0_49[11]), .sum(weight_1_49[7]), .cout(weight_1_50[6]));
full_adder fa291(.a(weight_0_50[8]), .b(weight_0_50[9]), .cin(weight_0_50[10]), .sum(weight_1_50[7]), .cout(weight_1_51[6]));
full_adder fa292(.a(weight_0_51[7]), .b(weight_0_51[8]), .cin(weight_0_51[9]), .sum(weight_1_51[7]), .cout(weight_1_52[4]));
full_adder fa293(.a(weight_0_52[6]), .b(weight_0_52[7]), .cin(weight_0_52[8]), .sum(weight_1_52[5]), .cout(weight_1_53[4]));
full_adder fa294(.a(weight_0_53[5]), .b(weight_0_53[6]), .cin(weight_0_53[7]), .sum(weight_1_53[5]), .cout(weight_1_54[4]));
full_adder fa295(.a(weight_0_54[4]), .b(weight_0_54[5]), .cin(weight_0_54[6]), .sum(weight_1_54[5]), .cout(weight_1_55[2]));
full_adder fa296(.a(weight_0_55[3]), .b(weight_0_55[4]), .cin(weight_0_55[5]), .sum(weight_1_55[3]), .cout(weight_1_56[2]));
full_adder fa297(.a(weight_0_56[2]), .b(weight_0_56[3]), .cin(weight_0_56[4]), .sum(weight_1_56[3]), .cout(weight_1_57[2]));
full_adder fa298(.a(weight_0_57[1]), .b(weight_0_57[2]), .cin(weight_0_57[3]), .sum(weight_1_57[3]), .cout(weight_1_58[0]));
full_adder fa299(.a(weight_0_58[0]), .b(weight_0_58[1]), .cin(weight_0_58[2]), .sum(weight_1_58[1]), .cout(weight_1_59[0]));
half_adder ha19(.a(weight_0_59[0]), .b(weight_0_59[1]), .sum(weight_1_59[1]), .cout(weight_1_60[0]));
assign weight_1_60[1] = weight_0_60[0];
assign weight_1_30[20] = weight_0_30[30];
assign weight_1_31[20] = weight_0_31[30];
assign weight_1_32[20] = weight_0_32[29];
assign weight_1_33[20] = weight_0_33[28];
assign weight_1_34[18] = weight_0_34[27];
assign weight_1_35[18] = weight_0_35[26];
assign weight_1_36[18] = weight_0_36[25];
assign weight_1_37[16] = weight_0_37[24];
assign weight_1_38[16] = weight_0_38[23];
assign weight_1_39[16] = weight_0_39[22];
assign weight_1_40[14] = weight_0_40[21];
assign weight_1_41[14] = weight_0_41[20];
assign weight_1_42[14] = weight_0_42[19];
assign weight_1_43[12] = weight_0_43[18];
assign weight_1_44[12] = weight_0_44[17];
assign weight_1_45[12] = weight_0_45[16];
assign weight_1_46[10] = weight_0_46[15];
assign weight_1_47[10] = weight_0_47[14];
assign weight_1_48[10] = weight_0_48[13];
assign weight_1_49[8] = weight_0_49[12];
assign weight_1_50[8] = weight_0_50[11];
assign weight_1_51[8] = weight_0_51[10];
assign weight_1_52[6] = weight_0_52[9];
assign weight_1_53[6] = weight_0_53[8];
assign weight_1_54[6] = weight_0_54[7];
assign weight_1_55[4] = weight_0_55[6];
assign weight_1_56[4] = weight_0_56[5];
assign weight_1_57[4] = weight_0_57[4];
assign weight_1_58[2] = weight_0_58[3];
assign weight_1_59[2] = weight_0_59[2];
assign weight_1_60[2] = weight_0_60[1];
assign weight_1_61[0] = weight_0_61[0];
assign weight_1_31[21] = weight_0_31[31];
assign weight_1_32[21] = weight_0_32[30];
assign weight_1_33[21] = weight_0_33[29];
assign weight_1_34[19] = weight_0_34[28];
assign weight_1_35[19] = weight_0_35[27];
assign weight_1_36[19] = weight_0_36[26];
assign weight_1_37[17] = weight_0_37[25];
assign weight_1_38[17] = weight_0_38[24];
assign weight_1_39[17] = weight_0_39[23];
assign weight_1_40[15] = weight_0_40[22];
assign weight_1_41[15] = weight_0_41[21];
assign weight_1_42[15] = weight_0_42[20];
assign weight_1_43[13] = weight_0_43[19];
assign weight_1_44[13] = weight_0_44[18];
assign weight_1_45[13] = weight_0_45[17];
assign weight_1_46[11] = weight_0_46[16];
assign weight_1_47[11] = weight_0_47[15];
assign weight_1_48[11] = weight_0_48[14];
assign weight_1_49[9] = weight_0_49[13];
assign weight_1_50[9] = weight_0_50[12];
assign weight_1_51[9] = weight_0_51[11];
assign weight_1_52[7] = weight_0_52[10];
assign weight_1_53[7] = weight_0_53[9];
assign weight_1_54[7] = weight_0_54[8];
assign weight_1_55[5] = weight_0_55[7];
assign weight_1_56[5] = weight_0_56[6];
assign weight_1_57[5] = weight_0_57[5];
assign weight_1_58[3] = weight_0_58[4];
assign weight_1_59[3] = weight_0_59[3];
assign weight_1_60[3] = weight_0_60[2];
assign weight_1_61[1] = weight_0_61[1];
assign weight_1_62 = weight_0_62;
logic weight_2_0;
logic weight_2_1;
logic weight_2_2;
logic [1:0] weight_2_3;
logic [1:0] weight_2_4;
logic [2:0] weight_2_5;
logic [2:0] weight_2_6;
logic [3:0] weight_2_7;
logic [3:0] weight_2_8;
logic [4:0] weight_2_9;
logic [4:0] weight_2_10;
logic [4:0] weight_2_11;
logic [5:0] weight_2_12;
logic [5:0] weight_2_13;
logic [6:0] weight_2_14;
logic [6:0] weight_2_15;
logic [7:0] weight_2_16;
logic [7:0] weight_2_17;
logic [8:0] weight_2_18;
logic [8:0] weight_2_19;
logic [8:0] weight_2_20;
logic [9:0] weight_2_21;
logic [9:0] weight_2_22;
logic [10:0] weight_2_23;
logic [10:0] weight_2_24;
logic [11:0] weight_2_25;
logic [11:0] weight_2_26;
logic [12:0] weight_2_27;
logic [12:0] weight_2_28;
logic [12:0] weight_2_29;
logic [13:0] weight_2_30;
logic [14:0] weight_2_31;
logic [14:0] weight_2_32;
logic [14:0] weight_2_33;
logic [14:0] weight_2_34;
logic [13:0] weight_2_35;
logic [13:0] weight_2_36;
logic [12:0] weight_2_37;
logic [12:0] weight_2_38;
logic [12:0] weight_2_39;
logic [11:0] weight_2_40;
logic [10:0] weight_2_41;
logic [10:0] weight_2_42;
logic [10:0] weight_2_43;
logic [9:0] weight_2_44;
logic [9:0] weight_2_45;
logic [8:0] weight_2_46;
logic [8:0] weight_2_47;
logic [8:0] weight_2_48;
logic [7:0] weight_2_49;
logic [6:0] weight_2_50;
logic [6:0] weight_2_51;
logic [6:0] weight_2_52;
logic [5:0] weight_2_53;
logic [5:0] weight_2_54;
logic [4:0] weight_2_55;
logic [4:0] weight_2_56;
logic [4:0] weight_2_57;
logic [3:0] weight_2_58;
logic [2:0] weight_2_59;
logic [2:0] weight_2_60;
logic [2:0] weight_2_61;
logic weight_2_62;

logic en_reg_1;
logic weight_2_0_reg;
logic weight_2_1_reg;
logic weight_2_2_reg;
logic [1:0] weight_2_3_reg;
logic [1:0] weight_2_4_reg;
logic [2:0] weight_2_5_reg;
logic [2:0] weight_2_6_reg;
logic [3:0] weight_2_7_reg;
logic [3:0] weight_2_8_reg;
logic [4:0] weight_2_9_reg;
logic [4:0] weight_2_10_reg;
logic [4:0] weight_2_11_reg;
logic [5:0] weight_2_12_reg;
logic [5:0] weight_2_13_reg;
logic [6:0] weight_2_14_reg;
logic [6:0] weight_2_15_reg;
logic [7:0] weight_2_16_reg;
logic [7:0] weight_2_17_reg;
logic [8:0] weight_2_18_reg;
logic [8:0] weight_2_19_reg;
logic [8:0] weight_2_20_reg;
logic [9:0] weight_2_21_reg;
logic [9:0] weight_2_22_reg;
logic [10:0] weight_2_23_reg;
logic [10:0] weight_2_24_reg;
logic [11:0] weight_2_25_reg;
logic [11:0] weight_2_26_reg;
logic [12:0] weight_2_27_reg;
logic [12:0] weight_2_28_reg;
logic [12:0] weight_2_29_reg;
logic [13:0] weight_2_30_reg;
logic [14:0] weight_2_31_reg;
logic [14:0] weight_2_32_reg;
logic [14:0] weight_2_33_reg;
logic [14:0] weight_2_34_reg;
logic [13:0] weight_2_35_reg;
logic [13:0] weight_2_36_reg;
logic [12:0] weight_2_37_reg;
logic [12:0] weight_2_38_reg;
logic [12:0] weight_2_39_reg;
logic [11:0] weight_2_40_reg;
logic [10:0] weight_2_41_reg;
logic [10:0] weight_2_42_reg;
logic [10:0] weight_2_43_reg;
logic [9:0] weight_2_44_reg;
logic [9:0] weight_2_45_reg;
logic [8:0] weight_2_46_reg;
logic [8:0] weight_2_47_reg;
logic [8:0] weight_2_48_reg;
logic [7:0] weight_2_49_reg;
logic [6:0] weight_2_50_reg;
logic [6:0] weight_2_51_reg;
logic [6:0] weight_2_52_reg;
logic [5:0] weight_2_53_reg;
logic [5:0] weight_2_54_reg;
logic [4:0] weight_2_55_reg;
logic [4:0] weight_2_56_reg;
logic [4:0] weight_2_57_reg;
logic [3:0] weight_2_58_reg;
logic [2:0] weight_2_59_reg;
logic [2:0] weight_2_60_reg;
logic [2:0] weight_2_61_reg;
logic weight_2_62_reg;

// First pipeline stage
always_ff @(posedge clk, negedge nrst) begin
    if (~nrst | multiplier_if.ready) begin
        en_reg_1 <= '0;
        weight_2_0_reg <= '0;
        weight_2_1_reg <= '0;
        weight_2_2_reg <= '0;
        weight_2_3_reg <= '0;
        weight_2_4_reg <= '0;
        weight_2_5_reg <= '0;
        weight_2_6_reg <= '0;
        weight_2_7_reg <= '0;
        weight_2_8_reg <= '0;
        weight_2_9_reg <= '0;
        weight_2_10_reg <= '0;
        weight_2_11_reg <= '0;
        weight_2_12_reg <= '0;
        weight_2_13_reg <= '0;
        weight_2_14_reg <= '0;
        weight_2_15_reg <= '0;
        weight_2_16_reg <= '0;
        weight_2_17_reg <= '0;
        weight_2_18_reg <= '0;
        weight_2_19_reg <= '0;
        weight_2_20_reg <= '0;
        weight_2_21_reg <= '0;
        weight_2_22_reg <= '0;
        weight_2_23_reg <= '0;
        weight_2_24_reg <= '0;
        weight_2_25_reg <= '0;
        weight_2_26_reg <= '0;
        weight_2_27_reg <= '0;
        weight_2_28_reg <= '0;
        weight_2_29_reg <= '0;
        weight_2_30_reg <= '0;
        weight_2_31_reg <= '0;
        weight_2_32_reg <= '0;
        weight_2_33_reg <= '0;
        weight_2_34_reg <= '0;
        weight_2_35_reg <= '0;
        weight_2_36_reg <= '0;
        weight_2_37_reg <= '0;
        weight_2_38_reg <= '0;
        weight_2_39_reg <= '0;
        weight_2_40_reg <= '0;
        weight_2_41_reg <= '0;
        weight_2_42_reg <= '0;
        weight_2_43_reg <= '0;
        weight_2_44_reg <= '0;
        weight_2_45_reg <= '0;
        weight_2_46_reg <= '0;
        weight_2_47_reg <= '0;
        weight_2_48_reg <= '0;
        weight_2_49_reg <= '0;
        weight_2_50_reg <= '0;
        weight_2_51_reg <= '0;
        weight_2_52_reg <= '0;
        weight_2_53_reg <= '0;
        weight_2_54_reg <= '0;
        weight_2_55_reg <= '0;
        weight_2_56_reg <= '0;
        weight_2_57_reg <= '0;
        weight_2_58_reg <= '0;
        weight_2_59_reg <= '0;
        weight_2_60_reg <= '0;
        weight_2_61_reg <= '0;
        weight_2_62_reg <= '0;
    end else begin
        en_reg_1 <= multiplier_if.en;
        weight_2_0_reg <= weight_2_0;
        weight_2_1_reg <= weight_2_1;
        weight_2_2_reg <= weight_2_2;
        weight_2_3_reg <= weight_2_3;
        weight_2_4_reg <= weight_2_4;
        weight_2_5_reg <= weight_2_5;
        weight_2_6_reg <= weight_2_6;
        weight_2_7_reg <= weight_2_7;
        weight_2_8_reg <= weight_2_8;
        weight_2_9_reg <= weight_2_9;
        weight_2_10_reg <= weight_2_10;
        weight_2_11_reg <= weight_2_11;
        weight_2_12_reg <= weight_2_12;
        weight_2_13_reg <= weight_2_13;
        weight_2_14_reg <= weight_2_14;
        weight_2_15_reg <= weight_2_15;
        weight_2_16_reg <= weight_2_16;
        weight_2_17_reg <= weight_2_17;
        weight_2_18_reg <= weight_2_18;
        weight_2_19_reg <= weight_2_19;
        weight_2_20_reg <= weight_2_20;
        weight_2_21_reg <= weight_2_21;
        weight_2_22_reg <= weight_2_22;
        weight_2_23_reg <= weight_2_23;
        weight_2_24_reg <= weight_2_24;
        weight_2_25_reg <= weight_2_25;
        weight_2_26_reg <= weight_2_26;
        weight_2_27_reg <= weight_2_27;
        weight_2_28_reg <= weight_2_28;
        weight_2_29_reg <= weight_2_29;
        weight_2_30_reg <= weight_2_30;
        weight_2_31_reg <= weight_2_31;
        weight_2_32_reg <= weight_2_32;
        weight_2_33_reg <= weight_2_33;
        weight_2_34_reg <= weight_2_34;
        weight_2_35_reg <= weight_2_35;
        weight_2_36_reg <= weight_2_36;
        weight_2_37_reg <= weight_2_37;
        weight_2_38_reg <= weight_2_38;
        weight_2_39_reg <= weight_2_39;
        weight_2_40_reg <= weight_2_40;
        weight_2_41_reg <= weight_2_41;
        weight_2_42_reg <= weight_2_42;
        weight_2_43_reg <= weight_2_43;
        weight_2_44_reg <= weight_2_44;
        weight_2_45_reg <= weight_2_45;
        weight_2_46_reg <= weight_2_46;
        weight_2_47_reg <= weight_2_47;
        weight_2_48_reg <= weight_2_48;
        weight_2_49_reg <= weight_2_49;
        weight_2_50_reg <= weight_2_50;
        weight_2_51_reg <= weight_2_51;
        weight_2_52_reg <= weight_2_52;
        weight_2_53_reg <= weight_2_53;
        weight_2_54_reg <= weight_2_54;
        weight_2_55_reg <= weight_2_55;
        weight_2_56_reg <= weight_2_56;
        weight_2_57_reg <= weight_2_57;
        weight_2_58_reg <= weight_2_58;
        weight_2_59_reg <= weight_2_59;
        weight_2_60_reg <= weight_2_60;
        weight_2_61_reg <= weight_2_61;
        weight_2_62_reg <= weight_2_62;
    end
end

assign weight_2_0 = weight_1_0;
assign weight_2_1 = weight_1_1;
half_adder ha20(.a(weight_1_2[0]), .b(weight_1_2[1]), .sum(weight_2_2), .cout(weight_2_3[0]));
full_adder fa300(.a(weight_1_3[0]), .b(weight_1_3[1]), .cin(weight_1_3[2]), .sum(weight_2_3[1]), .cout(weight_2_4[0]));
full_adder fa301(.a(weight_1_4[0]), .b(weight_1_4[1]), .cin(weight_1_4[2]), .sum(weight_2_4[1]), .cout(weight_2_5[0]));
full_adder fa302(.a(weight_1_5[0]), .b(weight_1_5[1]), .cin(weight_1_5[2]), .sum(weight_2_5[1]), .cout(weight_2_6[0]));
full_adder fa303(.a(weight_1_6[0]), .b(weight_1_6[1]), .cin(weight_1_6[2]), .sum(weight_2_6[1]), .cout(weight_2_7[0]));
full_adder fa304(.a(weight_1_7[0]), .b(weight_1_7[1]), .cin(weight_1_7[2]), .sum(weight_2_7[1]), .cout(weight_2_8[0]));
full_adder fa305(.a(weight_1_8[0]), .b(weight_1_8[1]), .cin(weight_1_8[2]), .sum(weight_2_8[1]), .cout(weight_2_9[0]));
full_adder fa306(.a(weight_1_9[0]), .b(weight_1_9[1]), .cin(weight_1_9[2]), .sum(weight_2_9[1]), .cout(weight_2_10[0]));
full_adder fa307(.a(weight_1_10[0]), .b(weight_1_10[1]), .cin(weight_1_10[2]), .sum(weight_2_10[1]), .cout(weight_2_11[0]));
full_adder fa308(.a(weight_1_11[0]), .b(weight_1_11[1]), .cin(weight_1_11[2]), .sum(weight_2_11[1]), .cout(weight_2_12[0]));
full_adder fa309(.a(weight_1_12[0]), .b(weight_1_12[1]), .cin(weight_1_12[2]), .sum(weight_2_12[1]), .cout(weight_2_13[0]));
full_adder fa310(.a(weight_1_13[0]), .b(weight_1_13[1]), .cin(weight_1_13[2]), .sum(weight_2_13[1]), .cout(weight_2_14[0]));
full_adder fa311(.a(weight_1_14[0]), .b(weight_1_14[1]), .cin(weight_1_14[2]), .sum(weight_2_14[1]), .cout(weight_2_15[0]));
full_adder fa312(.a(weight_1_15[0]), .b(weight_1_15[1]), .cin(weight_1_15[2]), .sum(weight_2_15[1]), .cout(weight_2_16[0]));
full_adder fa313(.a(weight_1_16[0]), .b(weight_1_16[1]), .cin(weight_1_16[2]), .sum(weight_2_16[1]), .cout(weight_2_17[0]));
full_adder fa314(.a(weight_1_17[0]), .b(weight_1_17[1]), .cin(weight_1_17[2]), .sum(weight_2_17[1]), .cout(weight_2_18[0]));
full_adder fa315(.a(weight_1_18[0]), .b(weight_1_18[1]), .cin(weight_1_18[2]), .sum(weight_2_18[1]), .cout(weight_2_19[0]));
full_adder fa316(.a(weight_1_19[0]), .b(weight_1_19[1]), .cin(weight_1_19[2]), .sum(weight_2_19[1]), .cout(weight_2_20[0]));
full_adder fa317(.a(weight_1_20[0]), .b(weight_1_20[1]), .cin(weight_1_20[2]), .sum(weight_2_20[1]), .cout(weight_2_21[0]));
full_adder fa318(.a(weight_1_21[0]), .b(weight_1_21[1]), .cin(weight_1_21[2]), .sum(weight_2_21[1]), .cout(weight_2_22[0]));
full_adder fa319(.a(weight_1_22[0]), .b(weight_1_22[1]), .cin(weight_1_22[2]), .sum(weight_2_22[1]), .cout(weight_2_23[0]));
full_adder fa320(.a(weight_1_23[0]), .b(weight_1_23[1]), .cin(weight_1_23[2]), .sum(weight_2_23[1]), .cout(weight_2_24[0]));
full_adder fa321(.a(weight_1_24[0]), .b(weight_1_24[1]), .cin(weight_1_24[2]), .sum(weight_2_24[1]), .cout(weight_2_25[0]));
full_adder fa322(.a(weight_1_25[0]), .b(weight_1_25[1]), .cin(weight_1_25[2]), .sum(weight_2_25[1]), .cout(weight_2_26[0]));
full_adder fa323(.a(weight_1_26[0]), .b(weight_1_26[1]), .cin(weight_1_26[2]), .sum(weight_2_26[1]), .cout(weight_2_27[0]));
full_adder fa324(.a(weight_1_27[0]), .b(weight_1_27[1]), .cin(weight_1_27[2]), .sum(weight_2_27[1]), .cout(weight_2_28[0]));
full_adder fa325(.a(weight_1_28[0]), .b(weight_1_28[1]), .cin(weight_1_28[2]), .sum(weight_2_28[1]), .cout(weight_2_29[0]));
full_adder fa326(.a(weight_1_29[0]), .b(weight_1_29[1]), .cin(weight_1_29[2]), .sum(weight_2_29[1]), .cout(weight_2_30[0]));
full_adder fa327(.a(weight_1_30[0]), .b(weight_1_30[1]), .cin(weight_1_30[2]), .sum(weight_2_30[1]), .cout(weight_2_31[0]));
full_adder fa328(.a(weight_1_31[0]), .b(weight_1_31[1]), .cin(weight_1_31[2]), .sum(weight_2_31[1]), .cout(weight_2_32[0]));
full_adder fa329(.a(weight_1_32[0]), .b(weight_1_32[1]), .cin(weight_1_32[2]), .sum(weight_2_32[1]), .cout(weight_2_33[0]));
full_adder fa330(.a(weight_1_33[0]), .b(weight_1_33[1]), .cin(weight_1_33[2]), .sum(weight_2_33[1]), .cout(weight_2_34[0]));
assign weight_2_34[1] = weight_1_34[0];
assign weight_2_35[0] = weight_1_35[0];
assign weight_2_36[0] = weight_1_36[0];
assign weight_2_5[2] = weight_1_5[3];
half_adder ha21(.a(weight_1_6[3]), .b(weight_1_6[4]), .sum(weight_2_6[2]), .cout(weight_2_7[2]));
half_adder ha22(.a(weight_1_7[3]), .b(weight_1_7[4]), .sum(weight_2_7[3]), .cout(weight_2_8[2]));
full_adder fa331(.a(weight_1_8[3]), .b(weight_1_8[4]), .cin(weight_1_8[5]), .sum(weight_2_8[3]), .cout(weight_2_9[2]));
full_adder fa332(.a(weight_1_9[3]), .b(weight_1_9[4]), .cin(weight_1_9[5]), .sum(weight_2_9[3]), .cout(weight_2_10[2]));
full_adder fa333(.a(weight_1_10[3]), .b(weight_1_10[4]), .cin(weight_1_10[5]), .sum(weight_2_10[3]), .cout(weight_2_11[2]));
full_adder fa334(.a(weight_1_11[3]), .b(weight_1_11[4]), .cin(weight_1_11[5]), .sum(weight_2_11[3]), .cout(weight_2_12[2]));
full_adder fa335(.a(weight_1_12[3]), .b(weight_1_12[4]), .cin(weight_1_12[5]), .sum(weight_2_12[3]), .cout(weight_2_13[2]));
full_adder fa336(.a(weight_1_13[3]), .b(weight_1_13[4]), .cin(weight_1_13[5]), .sum(weight_2_13[3]), .cout(weight_2_14[2]));
full_adder fa337(.a(weight_1_14[3]), .b(weight_1_14[4]), .cin(weight_1_14[5]), .sum(weight_2_14[3]), .cout(weight_2_15[2]));
full_adder fa338(.a(weight_1_15[3]), .b(weight_1_15[4]), .cin(weight_1_15[5]), .sum(weight_2_15[3]), .cout(weight_2_16[2]));
full_adder fa339(.a(weight_1_16[3]), .b(weight_1_16[4]), .cin(weight_1_16[5]), .sum(weight_2_16[3]), .cout(weight_2_17[2]));
full_adder fa340(.a(weight_1_17[3]), .b(weight_1_17[4]), .cin(weight_1_17[5]), .sum(weight_2_17[3]), .cout(weight_2_18[2]));
full_adder fa341(.a(weight_1_18[3]), .b(weight_1_18[4]), .cin(weight_1_18[5]), .sum(weight_2_18[3]), .cout(weight_2_19[2]));
full_adder fa342(.a(weight_1_19[3]), .b(weight_1_19[4]), .cin(weight_1_19[5]), .sum(weight_2_19[3]), .cout(weight_2_20[2]));
full_adder fa343(.a(weight_1_20[3]), .b(weight_1_20[4]), .cin(weight_1_20[5]), .sum(weight_2_20[3]), .cout(weight_2_21[2]));
full_adder fa344(.a(weight_1_21[3]), .b(weight_1_21[4]), .cin(weight_1_21[5]), .sum(weight_2_21[3]), .cout(weight_2_22[2]));
full_adder fa345(.a(weight_1_22[3]), .b(weight_1_22[4]), .cin(weight_1_22[5]), .sum(weight_2_22[3]), .cout(weight_2_23[2]));
full_adder fa346(.a(weight_1_23[3]), .b(weight_1_23[4]), .cin(weight_1_23[5]), .sum(weight_2_23[3]), .cout(weight_2_24[2]));
full_adder fa347(.a(weight_1_24[3]), .b(weight_1_24[4]), .cin(weight_1_24[5]), .sum(weight_2_24[3]), .cout(weight_2_25[2]));
full_adder fa348(.a(weight_1_25[3]), .b(weight_1_25[4]), .cin(weight_1_25[5]), .sum(weight_2_25[3]), .cout(weight_2_26[2]));
full_adder fa349(.a(weight_1_26[3]), .b(weight_1_26[4]), .cin(weight_1_26[5]), .sum(weight_2_26[3]), .cout(weight_2_27[2]));
full_adder fa350(.a(weight_1_27[3]), .b(weight_1_27[4]), .cin(weight_1_27[5]), .sum(weight_2_27[3]), .cout(weight_2_28[2]));
full_adder fa351(.a(weight_1_28[3]), .b(weight_1_28[4]), .cin(weight_1_28[5]), .sum(weight_2_28[3]), .cout(weight_2_29[2]));
full_adder fa352(.a(weight_1_29[3]), .b(weight_1_29[4]), .cin(weight_1_29[5]), .sum(weight_2_29[3]), .cout(weight_2_30[2]));
full_adder fa353(.a(weight_1_30[3]), .b(weight_1_30[4]), .cin(weight_1_30[5]), .sum(weight_2_30[3]), .cout(weight_2_31[2]));
full_adder fa354(.a(weight_1_31[3]), .b(weight_1_31[4]), .cin(weight_1_31[5]), .sum(weight_2_31[3]), .cout(weight_2_32[2]));
full_adder fa355(.a(weight_1_32[3]), .b(weight_1_32[4]), .cin(weight_1_32[5]), .sum(weight_2_32[3]), .cout(weight_2_33[2]));
full_adder fa356(.a(weight_1_33[3]), .b(weight_1_33[4]), .cin(weight_1_33[5]), .sum(weight_2_33[3]), .cout(weight_2_34[2]));
full_adder fa357(.a(weight_1_34[1]), .b(weight_1_34[2]), .cin(weight_1_34[3]), .sum(weight_2_34[3]), .cout(weight_2_35[1]));
full_adder fa358(.a(weight_1_35[1]), .b(weight_1_35[2]), .cin(weight_1_35[3]), .sum(weight_2_35[2]), .cout(weight_2_36[1]));
full_adder fa359(.a(weight_1_36[1]), .b(weight_1_36[2]), .cin(weight_1_36[3]), .sum(weight_2_36[2]), .cout(weight_2_37[0]));
half_adder ha23(.a(weight_1_37[0]), .b(weight_1_37[1]), .sum(weight_2_37[1]), .cout(weight_2_38[0]));
half_adder ha24(.a(weight_1_38[0]), .b(weight_1_38[1]), .sum(weight_2_38[1]), .cout(weight_2_39[0]));
half_adder ha25(.a(weight_1_39[0]), .b(weight_1_39[1]), .sum(weight_2_39[1]), .cout(weight_2_40[0]));
assign weight_2_9[4] = weight_1_9[6];
assign weight_2_10[4] = weight_1_10[6];
half_adder ha26(.a(weight_1_11[6]), .b(weight_1_11[7]), .sum(weight_2_11[4]), .cout(weight_2_12[4]));
full_adder fa360(.a(weight_1_12[6]), .b(weight_1_12[7]), .cin(weight_1_12[8]), .sum(weight_2_12[5]), .cout(weight_2_13[4]));
full_adder fa361(.a(weight_1_13[6]), .b(weight_1_13[7]), .cin(weight_1_13[8]), .sum(weight_2_13[5]), .cout(weight_2_14[4]));
full_adder fa362(.a(weight_1_14[6]), .b(weight_1_14[7]), .cin(weight_1_14[8]), .sum(weight_2_14[5]), .cout(weight_2_15[4]));
full_adder fa363(.a(weight_1_15[6]), .b(weight_1_15[7]), .cin(weight_1_15[8]), .sum(weight_2_15[5]), .cout(weight_2_16[4]));
full_adder fa364(.a(weight_1_16[6]), .b(weight_1_16[7]), .cin(weight_1_16[8]), .sum(weight_2_16[5]), .cout(weight_2_17[4]));
full_adder fa365(.a(weight_1_17[6]), .b(weight_1_17[7]), .cin(weight_1_17[8]), .sum(weight_2_17[5]), .cout(weight_2_18[4]));
full_adder fa366(.a(weight_1_18[6]), .b(weight_1_18[7]), .cin(weight_1_18[8]), .sum(weight_2_18[5]), .cout(weight_2_19[4]));
full_adder fa367(.a(weight_1_19[6]), .b(weight_1_19[7]), .cin(weight_1_19[8]), .sum(weight_2_19[5]), .cout(weight_2_20[4]));
full_adder fa368(.a(weight_1_20[6]), .b(weight_1_20[7]), .cin(weight_1_20[8]), .sum(weight_2_20[5]), .cout(weight_2_21[4]));
full_adder fa369(.a(weight_1_21[6]), .b(weight_1_21[7]), .cin(weight_1_21[8]), .sum(weight_2_21[5]), .cout(weight_2_22[4]));
full_adder fa370(.a(weight_1_22[6]), .b(weight_1_22[7]), .cin(weight_1_22[8]), .sum(weight_2_22[5]), .cout(weight_2_23[4]));
full_adder fa371(.a(weight_1_23[6]), .b(weight_1_23[7]), .cin(weight_1_23[8]), .sum(weight_2_23[5]), .cout(weight_2_24[4]));
full_adder fa372(.a(weight_1_24[6]), .b(weight_1_24[7]), .cin(weight_1_24[8]), .sum(weight_2_24[5]), .cout(weight_2_25[4]));
full_adder fa373(.a(weight_1_25[6]), .b(weight_1_25[7]), .cin(weight_1_25[8]), .sum(weight_2_25[5]), .cout(weight_2_26[4]));
full_adder fa374(.a(weight_1_26[6]), .b(weight_1_26[7]), .cin(weight_1_26[8]), .sum(weight_2_26[5]), .cout(weight_2_27[4]));
full_adder fa375(.a(weight_1_27[6]), .b(weight_1_27[7]), .cin(weight_1_27[8]), .sum(weight_2_27[5]), .cout(weight_2_28[4]));
full_adder fa376(.a(weight_1_28[6]), .b(weight_1_28[7]), .cin(weight_1_28[8]), .sum(weight_2_28[5]), .cout(weight_2_29[4]));
full_adder fa377(.a(weight_1_29[6]), .b(weight_1_29[7]), .cin(weight_1_29[8]), .sum(weight_2_29[5]), .cout(weight_2_30[4]));
full_adder fa378(.a(weight_1_30[6]), .b(weight_1_30[7]), .cin(weight_1_30[8]), .sum(weight_2_30[5]), .cout(weight_2_31[4]));
full_adder fa379(.a(weight_1_31[6]), .b(weight_1_31[7]), .cin(weight_1_31[8]), .sum(weight_2_31[5]), .cout(weight_2_32[4]));
full_adder fa380(.a(weight_1_32[6]), .b(weight_1_32[7]), .cin(weight_1_32[8]), .sum(weight_2_32[5]), .cout(weight_2_33[4]));
full_adder fa381(.a(weight_1_33[6]), .b(weight_1_33[7]), .cin(weight_1_33[8]), .sum(weight_2_33[5]), .cout(weight_2_34[4]));
full_adder fa382(.a(weight_1_34[4]), .b(weight_1_34[5]), .cin(weight_1_34[6]), .sum(weight_2_34[5]), .cout(weight_2_35[3]));
full_adder fa383(.a(weight_1_35[4]), .b(weight_1_35[5]), .cin(weight_1_35[6]), .sum(weight_2_35[4]), .cout(weight_2_36[3]));
full_adder fa384(.a(weight_1_36[4]), .b(weight_1_36[5]), .cin(weight_1_36[6]), .sum(weight_2_36[4]), .cout(weight_2_37[2]));
full_adder fa385(.a(weight_1_37[2]), .b(weight_1_37[3]), .cin(weight_1_37[4]), .sum(weight_2_37[3]), .cout(weight_2_38[2]));
full_adder fa386(.a(weight_1_38[2]), .b(weight_1_38[3]), .cin(weight_1_38[4]), .sum(weight_2_38[3]), .cout(weight_2_39[2]));
full_adder fa387(.a(weight_1_39[2]), .b(weight_1_39[3]), .cin(weight_1_39[4]), .sum(weight_2_39[3]), .cout(weight_2_40[1]));
full_adder fa388(.a(weight_1_40[0]), .b(weight_1_40[1]), .cin(weight_1_40[2]), .sum(weight_2_40[2]), .cout(weight_2_41[0]));
full_adder fa389(.a(weight_1_41[0]), .b(weight_1_41[1]), .cin(weight_1_41[2]), .sum(weight_2_41[1]), .cout(weight_2_42[0]));
full_adder fa390(.a(weight_1_42[0]), .b(weight_1_42[1]), .cin(weight_1_42[2]), .sum(weight_2_42[1]), .cout(weight_2_43[0]));
assign weight_2_43[1] = weight_1_43[0];
assign weight_2_44[0] = weight_1_44[0];
assign weight_2_45[0] = weight_1_45[0];
assign weight_2_14[6] = weight_1_14[9];
half_adder ha27(.a(weight_1_15[9]), .b(weight_1_15[10]), .sum(weight_2_15[6]), .cout(weight_2_16[6]));
half_adder ha28(.a(weight_1_16[9]), .b(weight_1_16[10]), .sum(weight_2_16[7]), .cout(weight_2_17[6]));
full_adder fa391(.a(weight_1_17[9]), .b(weight_1_17[10]), .cin(weight_1_17[11]), .sum(weight_2_17[7]), .cout(weight_2_18[6]));
full_adder fa392(.a(weight_1_18[9]), .b(weight_1_18[10]), .cin(weight_1_18[11]), .sum(weight_2_18[7]), .cout(weight_2_19[6]));
full_adder fa393(.a(weight_1_19[9]), .b(weight_1_19[10]), .cin(weight_1_19[11]), .sum(weight_2_19[7]), .cout(weight_2_20[6]));
full_adder fa394(.a(weight_1_20[9]), .b(weight_1_20[10]), .cin(weight_1_20[11]), .sum(weight_2_20[7]), .cout(weight_2_21[6]));
full_adder fa395(.a(weight_1_21[9]), .b(weight_1_21[10]), .cin(weight_1_21[11]), .sum(weight_2_21[7]), .cout(weight_2_22[6]));
full_adder fa396(.a(weight_1_22[9]), .b(weight_1_22[10]), .cin(weight_1_22[11]), .sum(weight_2_22[7]), .cout(weight_2_23[6]));
full_adder fa397(.a(weight_1_23[9]), .b(weight_1_23[10]), .cin(weight_1_23[11]), .sum(weight_2_23[7]), .cout(weight_2_24[6]));
full_adder fa398(.a(weight_1_24[9]), .b(weight_1_24[10]), .cin(weight_1_24[11]), .sum(weight_2_24[7]), .cout(weight_2_25[6]));
full_adder fa399(.a(weight_1_25[9]), .b(weight_1_25[10]), .cin(weight_1_25[11]), .sum(weight_2_25[7]), .cout(weight_2_26[6]));
full_adder fa400(.a(weight_1_26[9]), .b(weight_1_26[10]), .cin(weight_1_26[11]), .sum(weight_2_26[7]), .cout(weight_2_27[6]));
full_adder fa401(.a(weight_1_27[9]), .b(weight_1_27[10]), .cin(weight_1_27[11]), .sum(weight_2_27[7]), .cout(weight_2_28[6]));
full_adder fa402(.a(weight_1_28[9]), .b(weight_1_28[10]), .cin(weight_1_28[11]), .sum(weight_2_28[7]), .cout(weight_2_29[6]));
full_adder fa403(.a(weight_1_29[9]), .b(weight_1_29[10]), .cin(weight_1_29[11]), .sum(weight_2_29[7]), .cout(weight_2_30[6]));
full_adder fa404(.a(weight_1_30[9]), .b(weight_1_30[10]), .cin(weight_1_30[11]), .sum(weight_2_30[7]), .cout(weight_2_31[6]));
full_adder fa405(.a(weight_1_31[9]), .b(weight_1_31[10]), .cin(weight_1_31[11]), .sum(weight_2_31[7]), .cout(weight_2_32[6]));
full_adder fa406(.a(weight_1_32[9]), .b(weight_1_32[10]), .cin(weight_1_32[11]), .sum(weight_2_32[7]), .cout(weight_2_33[6]));
full_adder fa407(.a(weight_1_33[9]), .b(weight_1_33[10]), .cin(weight_1_33[11]), .sum(weight_2_33[7]), .cout(weight_2_34[6]));
full_adder fa408(.a(weight_1_34[7]), .b(weight_1_34[8]), .cin(weight_1_34[9]), .sum(weight_2_34[7]), .cout(weight_2_35[5]));
full_adder fa409(.a(weight_1_35[7]), .b(weight_1_35[8]), .cin(weight_1_35[9]), .sum(weight_2_35[6]), .cout(weight_2_36[5]));
full_adder fa410(.a(weight_1_36[7]), .b(weight_1_36[8]), .cin(weight_1_36[9]), .sum(weight_2_36[6]), .cout(weight_2_37[4]));
full_adder fa411(.a(weight_1_37[5]), .b(weight_1_37[6]), .cin(weight_1_37[7]), .sum(weight_2_37[5]), .cout(weight_2_38[4]));
full_adder fa412(.a(weight_1_38[5]), .b(weight_1_38[6]), .cin(weight_1_38[7]), .sum(weight_2_38[5]), .cout(weight_2_39[4]));
full_adder fa413(.a(weight_1_39[5]), .b(weight_1_39[6]), .cin(weight_1_39[7]), .sum(weight_2_39[5]), .cout(weight_2_40[3]));
full_adder fa414(.a(weight_1_40[3]), .b(weight_1_40[4]), .cin(weight_1_40[5]), .sum(weight_2_40[4]), .cout(weight_2_41[2]));
full_adder fa415(.a(weight_1_41[3]), .b(weight_1_41[4]), .cin(weight_1_41[5]), .sum(weight_2_41[3]), .cout(weight_2_42[2]));
full_adder fa416(.a(weight_1_42[3]), .b(weight_1_42[4]), .cin(weight_1_42[5]), .sum(weight_2_42[3]), .cout(weight_2_43[2]));
full_adder fa417(.a(weight_1_43[1]), .b(weight_1_43[2]), .cin(weight_1_43[3]), .sum(weight_2_43[3]), .cout(weight_2_44[1]));
full_adder fa418(.a(weight_1_44[1]), .b(weight_1_44[2]), .cin(weight_1_44[3]), .sum(weight_2_44[2]), .cout(weight_2_45[1]));
full_adder fa419(.a(weight_1_45[1]), .b(weight_1_45[2]), .cin(weight_1_45[3]), .sum(weight_2_45[2]), .cout(weight_2_46[0]));
half_adder ha29(.a(weight_1_46[0]), .b(weight_1_46[1]), .sum(weight_2_46[1]), .cout(weight_2_47[0]));
half_adder ha30(.a(weight_1_47[0]), .b(weight_1_47[1]), .sum(weight_2_47[1]), .cout(weight_2_48[0]));
half_adder ha31(.a(weight_1_48[0]), .b(weight_1_48[1]), .sum(weight_2_48[1]), .cout(weight_2_49[0]));
assign weight_2_18[8] = weight_1_18[12];
assign weight_2_19[8] = weight_1_19[12];
half_adder ha32(.a(weight_1_20[12]), .b(weight_1_20[13]), .sum(weight_2_20[8]), .cout(weight_2_21[8]));
full_adder fa420(.a(weight_1_21[12]), .b(weight_1_21[13]), .cin(weight_1_21[14]), .sum(weight_2_21[9]), .cout(weight_2_22[8]));
full_adder fa421(.a(weight_1_22[12]), .b(weight_1_22[13]), .cin(weight_1_22[14]), .sum(weight_2_22[9]), .cout(weight_2_23[8]));
full_adder fa422(.a(weight_1_23[12]), .b(weight_1_23[13]), .cin(weight_1_23[14]), .sum(weight_2_23[9]), .cout(weight_2_24[8]));
full_adder fa423(.a(weight_1_24[12]), .b(weight_1_24[13]), .cin(weight_1_24[14]), .sum(weight_2_24[9]), .cout(weight_2_25[8]));
full_adder fa424(.a(weight_1_25[12]), .b(weight_1_25[13]), .cin(weight_1_25[14]), .sum(weight_2_25[9]), .cout(weight_2_26[8]));
full_adder fa425(.a(weight_1_26[12]), .b(weight_1_26[13]), .cin(weight_1_26[14]), .sum(weight_2_26[9]), .cout(weight_2_27[8]));
full_adder fa426(.a(weight_1_27[12]), .b(weight_1_27[13]), .cin(weight_1_27[14]), .sum(weight_2_27[9]), .cout(weight_2_28[8]));
full_adder fa427(.a(weight_1_28[12]), .b(weight_1_28[13]), .cin(weight_1_28[14]), .sum(weight_2_28[9]), .cout(weight_2_29[8]));
full_adder fa428(.a(weight_1_29[12]), .b(weight_1_29[13]), .cin(weight_1_29[14]), .sum(weight_2_29[9]), .cout(weight_2_30[8]));
full_adder fa429(.a(weight_1_30[12]), .b(weight_1_30[13]), .cin(weight_1_30[14]), .sum(weight_2_30[9]), .cout(weight_2_31[8]));
full_adder fa430(.a(weight_1_31[12]), .b(weight_1_31[13]), .cin(weight_1_31[14]), .sum(weight_2_31[9]), .cout(weight_2_32[8]));
full_adder fa431(.a(weight_1_32[12]), .b(weight_1_32[13]), .cin(weight_1_32[14]), .sum(weight_2_32[9]), .cout(weight_2_33[8]));
full_adder fa432(.a(weight_1_33[12]), .b(weight_1_33[13]), .cin(weight_1_33[14]), .sum(weight_2_33[9]), .cout(weight_2_34[8]));
full_adder fa433(.a(weight_1_34[10]), .b(weight_1_34[11]), .cin(weight_1_34[12]), .sum(weight_2_34[9]), .cout(weight_2_35[7]));
full_adder fa434(.a(weight_1_35[10]), .b(weight_1_35[11]), .cin(weight_1_35[12]), .sum(weight_2_35[8]), .cout(weight_2_36[7]));
full_adder fa435(.a(weight_1_36[10]), .b(weight_1_36[11]), .cin(weight_1_36[12]), .sum(weight_2_36[8]), .cout(weight_2_37[6]));
full_adder fa436(.a(weight_1_37[8]), .b(weight_1_37[9]), .cin(weight_1_37[10]), .sum(weight_2_37[7]), .cout(weight_2_38[6]));
full_adder fa437(.a(weight_1_38[8]), .b(weight_1_38[9]), .cin(weight_1_38[10]), .sum(weight_2_38[7]), .cout(weight_2_39[6]));
full_adder fa438(.a(weight_1_39[8]), .b(weight_1_39[9]), .cin(weight_1_39[10]), .sum(weight_2_39[7]), .cout(weight_2_40[5]));
full_adder fa439(.a(weight_1_40[6]), .b(weight_1_40[7]), .cin(weight_1_40[8]), .sum(weight_2_40[6]), .cout(weight_2_41[4]));
full_adder fa440(.a(weight_1_41[6]), .b(weight_1_41[7]), .cin(weight_1_41[8]), .sum(weight_2_41[5]), .cout(weight_2_42[4]));
full_adder fa441(.a(weight_1_42[6]), .b(weight_1_42[7]), .cin(weight_1_42[8]), .sum(weight_2_42[5]), .cout(weight_2_43[4]));
full_adder fa442(.a(weight_1_43[4]), .b(weight_1_43[5]), .cin(weight_1_43[6]), .sum(weight_2_43[5]), .cout(weight_2_44[3]));
full_adder fa443(.a(weight_1_44[4]), .b(weight_1_44[5]), .cin(weight_1_44[6]), .sum(weight_2_44[4]), .cout(weight_2_45[3]));
full_adder fa444(.a(weight_1_45[4]), .b(weight_1_45[5]), .cin(weight_1_45[6]), .sum(weight_2_45[4]), .cout(weight_2_46[2]));
full_adder fa445(.a(weight_1_46[2]), .b(weight_1_46[3]), .cin(weight_1_46[4]), .sum(weight_2_46[3]), .cout(weight_2_47[2]));
full_adder fa446(.a(weight_1_47[2]), .b(weight_1_47[3]), .cin(weight_1_47[4]), .sum(weight_2_47[3]), .cout(weight_2_48[2]));
full_adder fa447(.a(weight_1_48[2]), .b(weight_1_48[3]), .cin(weight_1_48[4]), .sum(weight_2_48[3]), .cout(weight_2_49[1]));
full_adder fa448(.a(weight_1_49[0]), .b(weight_1_49[1]), .cin(weight_1_49[2]), .sum(weight_2_49[2]), .cout(weight_2_50[0]));
full_adder fa449(.a(weight_1_50[0]), .b(weight_1_50[1]), .cin(weight_1_50[2]), .sum(weight_2_50[1]), .cout(weight_2_51[0]));
full_adder fa450(.a(weight_1_51[0]), .b(weight_1_51[1]), .cin(weight_1_51[2]), .sum(weight_2_51[1]), .cout(weight_2_52[0]));
assign weight_2_52[1] = weight_1_52[0];
assign weight_2_53[0] = weight_1_53[0];
assign weight_2_54[0] = weight_1_54[0];
assign weight_2_23[10] = weight_1_23[15];
half_adder ha33(.a(weight_1_24[15]), .b(weight_1_24[16]), .sum(weight_2_24[10]), .cout(weight_2_25[10]));
half_adder ha34(.a(weight_1_25[15]), .b(weight_1_25[16]), .sum(weight_2_25[11]), .cout(weight_2_26[10]));
full_adder fa451(.a(weight_1_26[15]), .b(weight_1_26[16]), .cin(weight_1_26[17]), .sum(weight_2_26[11]), .cout(weight_2_27[10]));
full_adder fa452(.a(weight_1_27[15]), .b(weight_1_27[16]), .cin(weight_1_27[17]), .sum(weight_2_27[11]), .cout(weight_2_28[10]));
full_adder fa453(.a(weight_1_28[15]), .b(weight_1_28[16]), .cin(weight_1_28[17]), .sum(weight_2_28[11]), .cout(weight_2_29[10]));
full_adder fa454(.a(weight_1_29[15]), .b(weight_1_29[16]), .cin(weight_1_29[17]), .sum(weight_2_29[11]), .cout(weight_2_30[10]));
full_adder fa455(.a(weight_1_30[15]), .b(weight_1_30[16]), .cin(weight_1_30[17]), .sum(weight_2_30[11]), .cout(weight_2_31[10]));
full_adder fa456(.a(weight_1_31[15]), .b(weight_1_31[16]), .cin(weight_1_31[17]), .sum(weight_2_31[11]), .cout(weight_2_32[10]));
full_adder fa457(.a(weight_1_32[15]), .b(weight_1_32[16]), .cin(weight_1_32[17]), .sum(weight_2_32[11]), .cout(weight_2_33[10]));
full_adder fa458(.a(weight_1_33[15]), .b(weight_1_33[16]), .cin(weight_1_33[17]), .sum(weight_2_33[11]), .cout(weight_2_34[10]));
full_adder fa459(.a(weight_1_34[13]), .b(weight_1_34[14]), .cin(weight_1_34[15]), .sum(weight_2_34[11]), .cout(weight_2_35[9]));
full_adder fa460(.a(weight_1_35[13]), .b(weight_1_35[14]), .cin(weight_1_35[15]), .sum(weight_2_35[10]), .cout(weight_2_36[9]));
full_adder fa461(.a(weight_1_36[13]), .b(weight_1_36[14]), .cin(weight_1_36[15]), .sum(weight_2_36[10]), .cout(weight_2_37[8]));
full_adder fa462(.a(weight_1_37[11]), .b(weight_1_37[12]), .cin(weight_1_37[13]), .sum(weight_2_37[9]), .cout(weight_2_38[8]));
full_adder fa463(.a(weight_1_38[11]), .b(weight_1_38[12]), .cin(weight_1_38[13]), .sum(weight_2_38[9]), .cout(weight_2_39[8]));
full_adder fa464(.a(weight_1_39[11]), .b(weight_1_39[12]), .cin(weight_1_39[13]), .sum(weight_2_39[9]), .cout(weight_2_40[7]));
full_adder fa465(.a(weight_1_40[9]), .b(weight_1_40[10]), .cin(weight_1_40[11]), .sum(weight_2_40[8]), .cout(weight_2_41[6]));
full_adder fa466(.a(weight_1_41[9]), .b(weight_1_41[10]), .cin(weight_1_41[11]), .sum(weight_2_41[7]), .cout(weight_2_42[6]));
full_adder fa467(.a(weight_1_42[9]), .b(weight_1_42[10]), .cin(weight_1_42[11]), .sum(weight_2_42[7]), .cout(weight_2_43[6]));
full_adder fa468(.a(weight_1_43[7]), .b(weight_1_43[8]), .cin(weight_1_43[9]), .sum(weight_2_43[7]), .cout(weight_2_44[5]));
full_adder fa469(.a(weight_1_44[7]), .b(weight_1_44[8]), .cin(weight_1_44[9]), .sum(weight_2_44[6]), .cout(weight_2_45[5]));
full_adder fa470(.a(weight_1_45[7]), .b(weight_1_45[8]), .cin(weight_1_45[9]), .sum(weight_2_45[6]), .cout(weight_2_46[4]));
full_adder fa471(.a(weight_1_46[5]), .b(weight_1_46[6]), .cin(weight_1_46[7]), .sum(weight_2_46[5]), .cout(weight_2_47[4]));
full_adder fa472(.a(weight_1_47[5]), .b(weight_1_47[6]), .cin(weight_1_47[7]), .sum(weight_2_47[5]), .cout(weight_2_48[4]));
full_adder fa473(.a(weight_1_48[5]), .b(weight_1_48[6]), .cin(weight_1_48[7]), .sum(weight_2_48[5]), .cout(weight_2_49[3]));
full_adder fa474(.a(weight_1_49[3]), .b(weight_1_49[4]), .cin(weight_1_49[5]), .sum(weight_2_49[4]), .cout(weight_2_50[2]));
full_adder fa475(.a(weight_1_50[3]), .b(weight_1_50[4]), .cin(weight_1_50[5]), .sum(weight_2_50[3]), .cout(weight_2_51[2]));
full_adder fa476(.a(weight_1_51[3]), .b(weight_1_51[4]), .cin(weight_1_51[5]), .sum(weight_2_51[3]), .cout(weight_2_52[2]));
full_adder fa477(.a(weight_1_52[1]), .b(weight_1_52[2]), .cin(weight_1_52[3]), .sum(weight_2_52[3]), .cout(weight_2_53[1]));
full_adder fa478(.a(weight_1_53[1]), .b(weight_1_53[2]), .cin(weight_1_53[3]), .sum(weight_2_53[2]), .cout(weight_2_54[1]));
full_adder fa479(.a(weight_1_54[1]), .b(weight_1_54[2]), .cin(weight_1_54[3]), .sum(weight_2_54[2]), .cout(weight_2_55[0]));
half_adder ha35(.a(weight_1_55[0]), .b(weight_1_55[1]), .sum(weight_2_55[1]), .cout(weight_2_56[0]));
half_adder ha36(.a(weight_1_56[0]), .b(weight_1_56[1]), .sum(weight_2_56[1]), .cout(weight_2_57[0]));
half_adder ha37(.a(weight_1_57[0]), .b(weight_1_57[1]), .sum(weight_2_57[1]), .cout(weight_2_58[0]));
assign weight_2_27[12] = weight_1_27[18];
assign weight_2_28[12] = weight_1_28[18];
half_adder ha38(.a(weight_1_29[18]), .b(weight_1_29[19]), .sum(weight_2_29[12]), .cout(weight_2_30[12]));
full_adder fa480(.a(weight_1_30[18]), .b(weight_1_30[19]), .cin(weight_1_30[20]), .sum(weight_2_30[13]), .cout(weight_2_31[12]));
full_adder fa481(.a(weight_1_31[18]), .b(weight_1_31[19]), .cin(weight_1_31[20]), .sum(weight_2_31[13]), .cout(weight_2_32[12]));
full_adder fa482(.a(weight_1_32[18]), .b(weight_1_32[19]), .cin(weight_1_32[20]), .sum(weight_2_32[13]), .cout(weight_2_33[12]));
full_adder fa483(.a(weight_1_33[18]), .b(weight_1_33[19]), .cin(weight_1_33[20]), .sum(weight_2_33[13]), .cout(weight_2_34[12]));
full_adder fa484(.a(weight_1_34[16]), .b(weight_1_34[17]), .cin(weight_1_34[18]), .sum(weight_2_34[13]), .cout(weight_2_35[11]));
full_adder fa485(.a(weight_1_35[16]), .b(weight_1_35[17]), .cin(weight_1_35[18]), .sum(weight_2_35[12]), .cout(weight_2_36[11]));
full_adder fa486(.a(weight_1_36[16]), .b(weight_1_36[17]), .cin(weight_1_36[18]), .sum(weight_2_36[12]), .cout(weight_2_37[10]));
full_adder fa487(.a(weight_1_37[14]), .b(weight_1_37[15]), .cin(weight_1_37[16]), .sum(weight_2_37[11]), .cout(weight_2_38[10]));
full_adder fa488(.a(weight_1_38[14]), .b(weight_1_38[15]), .cin(weight_1_38[16]), .sum(weight_2_38[11]), .cout(weight_2_39[10]));
full_adder fa489(.a(weight_1_39[14]), .b(weight_1_39[15]), .cin(weight_1_39[16]), .sum(weight_2_39[11]), .cout(weight_2_40[9]));
full_adder fa490(.a(weight_1_40[12]), .b(weight_1_40[13]), .cin(weight_1_40[14]), .sum(weight_2_40[10]), .cout(weight_2_41[8]));
full_adder fa491(.a(weight_1_41[12]), .b(weight_1_41[13]), .cin(weight_1_41[14]), .sum(weight_2_41[9]), .cout(weight_2_42[8]));
full_adder fa492(.a(weight_1_42[12]), .b(weight_1_42[13]), .cin(weight_1_42[14]), .sum(weight_2_42[9]), .cout(weight_2_43[8]));
full_adder fa493(.a(weight_1_43[10]), .b(weight_1_43[11]), .cin(weight_1_43[12]), .sum(weight_2_43[9]), .cout(weight_2_44[7]));
full_adder fa494(.a(weight_1_44[10]), .b(weight_1_44[11]), .cin(weight_1_44[12]), .sum(weight_2_44[8]), .cout(weight_2_45[7]));
full_adder fa495(.a(weight_1_45[10]), .b(weight_1_45[11]), .cin(weight_1_45[12]), .sum(weight_2_45[8]), .cout(weight_2_46[6]));
full_adder fa496(.a(weight_1_46[8]), .b(weight_1_46[9]), .cin(weight_1_46[10]), .sum(weight_2_46[7]), .cout(weight_2_47[6]));
full_adder fa497(.a(weight_1_47[8]), .b(weight_1_47[9]), .cin(weight_1_47[10]), .sum(weight_2_47[7]), .cout(weight_2_48[6]));
full_adder fa498(.a(weight_1_48[8]), .b(weight_1_48[9]), .cin(weight_1_48[10]), .sum(weight_2_48[7]), .cout(weight_2_49[5]));
full_adder fa499(.a(weight_1_49[6]), .b(weight_1_49[7]), .cin(weight_1_49[8]), .sum(weight_2_49[6]), .cout(weight_2_50[4]));
full_adder fa500(.a(weight_1_50[6]), .b(weight_1_50[7]), .cin(weight_1_50[8]), .sum(weight_2_50[5]), .cout(weight_2_51[4]));
full_adder fa501(.a(weight_1_51[6]), .b(weight_1_51[7]), .cin(weight_1_51[8]), .sum(weight_2_51[5]), .cout(weight_2_52[4]));
full_adder fa502(.a(weight_1_52[4]), .b(weight_1_52[5]), .cin(weight_1_52[6]), .sum(weight_2_52[5]), .cout(weight_2_53[3]));
full_adder fa503(.a(weight_1_53[4]), .b(weight_1_53[5]), .cin(weight_1_53[6]), .sum(weight_2_53[4]), .cout(weight_2_54[3]));
full_adder fa504(.a(weight_1_54[4]), .b(weight_1_54[5]), .cin(weight_1_54[6]), .sum(weight_2_54[4]), .cout(weight_2_55[2]));
full_adder fa505(.a(weight_1_55[2]), .b(weight_1_55[3]), .cin(weight_1_55[4]), .sum(weight_2_55[3]), .cout(weight_2_56[2]));
full_adder fa506(.a(weight_1_56[2]), .b(weight_1_56[3]), .cin(weight_1_56[4]), .sum(weight_2_56[3]), .cout(weight_2_57[2]));
full_adder fa507(.a(weight_1_57[2]), .b(weight_1_57[3]), .cin(weight_1_57[4]), .sum(weight_2_57[3]), .cout(weight_2_58[1]));
full_adder fa508(.a(weight_1_58[0]), .b(weight_1_58[1]), .cin(weight_1_58[2]), .sum(weight_2_58[2]), .cout(weight_2_59[0]));
full_adder fa509(.a(weight_1_59[0]), .b(weight_1_59[1]), .cin(weight_1_59[2]), .sum(weight_2_59[1]), .cout(weight_2_60[0]));
full_adder fa510(.a(weight_1_60[0]), .b(weight_1_60[1]), .cin(weight_1_60[2]), .sum(weight_2_60[1]), .cout(weight_2_61[0]));
assign weight_2_61[1] = weight_1_61[0];
assign weight_2_31[14] = weight_1_31[21];
assign weight_2_32[14] = weight_1_32[21];
assign weight_2_33[14] = weight_1_33[21];
assign weight_2_34[14] = weight_1_34[19];
assign weight_2_35[13] = weight_1_35[19];
assign weight_2_36[13] = weight_1_36[19];
assign weight_2_37[12] = weight_1_37[17];
assign weight_2_38[12] = weight_1_38[17];
assign weight_2_39[12] = weight_1_39[17];
assign weight_2_40[11] = weight_1_40[15];
assign weight_2_41[10] = weight_1_41[15];
assign weight_2_42[10] = weight_1_42[15];
assign weight_2_43[10] = weight_1_43[13];
assign weight_2_44[9] = weight_1_44[13];
assign weight_2_45[9] = weight_1_45[13];
assign weight_2_46[8] = weight_1_46[11];
assign weight_2_47[8] = weight_1_47[11];
assign weight_2_48[8] = weight_1_48[11];
assign weight_2_49[7] = weight_1_49[9];
assign weight_2_50[6] = weight_1_50[9];
assign weight_2_51[6] = weight_1_51[9];
assign weight_2_52[6] = weight_1_52[7];
assign weight_2_53[5] = weight_1_53[7];
assign weight_2_54[5] = weight_1_54[7];
assign weight_2_55[4] = weight_1_55[5];
assign weight_2_56[4] = weight_1_56[5];
assign weight_2_57[4] = weight_1_57[5];
assign weight_2_58[3] = weight_1_58[3];
assign weight_2_59[2] = weight_1_59[3];
assign weight_2_60[2] = weight_1_60[3];
assign weight_2_61[2] = weight_1_61[1];
assign weight_2_62 = weight_1_62;
logic weight_3_0;
logic weight_3_1;
logic weight_3_2;
logic weight_3_3;
logic [1:0] weight_3_4;
logic [1:0] weight_3_5;
logic [1:0] weight_3_6;
logic [2:0] weight_3_7;
logic [2:0] weight_3_8;
logic [2:0] weight_3_9;
logic [3:0] weight_3_10;
logic [3:0] weight_3_11;
logic [3:0] weight_3_12;
logic [3:0] weight_3_13;
logic [4:0] weight_3_14;
logic [4:0] weight_3_15;
logic [4:0] weight_3_16;
logic [5:0] weight_3_17;
logic [5:0] weight_3_18;
logic [5:0] weight_3_19;
logic [5:0] weight_3_20;
logic [6:0] weight_3_21;
logic [6:0] weight_3_22;
logic [6:0] weight_3_23;
logic [7:0] weight_3_24;
logic [7:0] weight_3_25;
logic [7:0] weight_3_26;
logic [8:0] weight_3_27;
logic [8:0] weight_3_28;
logic [8:0] weight_3_29;
logic [8:0] weight_3_30;
logic [9:0] weight_3_31;
logic [9:0] weight_3_32;
logic [9:0] weight_3_33;
logic [9:0] weight_3_34;
logic [9:0] weight_3_35;
logic [9:0] weight_3_36;
logic [9:0] weight_3_37;
logic [8:0] weight_3_38;
logic [8:0] weight_3_39;
logic [7:0] weight_3_40;
logic [7:0] weight_3_41;
logic [7:0] weight_3_42;
logic [7:0] weight_3_43;
logic [7:0] weight_3_44;
logic [6:0] weight_3_45;
logic [5:0] weight_3_46;
logic [5:0] weight_3_47;
logic [5:0] weight_3_48;
logic [5:0] weight_3_49;
logic [5:0] weight_3_50;
logic [4:0] weight_3_51;
logic [4:0] weight_3_52;
logic [3:0] weight_3_53;
logic [3:0] weight_3_54;
logic [3:0] weight_3_55;
logic [3:0] weight_3_56;
logic [3:0] weight_3_57;
logic [3:0] weight_3_58;
logic [1:0] weight_3_59;
logic [1:0] weight_3_60;
logic [1:0] weight_3_61;
logic [1:0] weight_3_62;
assign weight_3_0 = weight_2_0_reg;
assign weight_3_1 = weight_2_1_reg;
assign weight_3_2 = weight_2_2_reg;
half_adder ha39(.a(weight_2_3_reg[0]), .b(weight_2_3_reg[1]), .sum(weight_3_3), .cout(weight_3_4[0]));
half_adder ha40(.a(weight_2_4_reg[0]), .b(weight_2_4_reg[1]), .sum(weight_3_4[1]), .cout(weight_3_5[0]));
full_adder fa511(.a(weight_2_5_reg[0]), .b(weight_2_5_reg[1]), .cin(weight_2_5_reg[2]), .sum(weight_3_5[1]), .cout(weight_3_6[0]));
full_adder fa512(.a(weight_2_6_reg[0]), .b(weight_2_6_reg[1]), .cin(weight_2_6_reg[2]), .sum(weight_3_6[1]), .cout(weight_3_7[0]));
full_adder fa513(.a(weight_2_7_reg[0]), .b(weight_2_7_reg[1]), .cin(weight_2_7_reg[2]), .sum(weight_3_7[1]), .cout(weight_3_8[0]));
full_adder fa514(.a(weight_2_8_reg[0]), .b(weight_2_8_reg[1]), .cin(weight_2_8_reg[2]), .sum(weight_3_8[1]), .cout(weight_3_9[0]));
full_adder fa515(.a(weight_2_9_reg[0]), .b(weight_2_9_reg[1]), .cin(weight_2_9_reg[2]), .sum(weight_3_9[1]), .cout(weight_3_10[0]));
full_adder fa516(.a(weight_2_10_reg[0]), .b(weight_2_10_reg[1]), .cin(weight_2_10_reg[2]), .sum(weight_3_10[1]), .cout(weight_3_11[0]));
full_adder fa517(.a(weight_2_11_reg[0]), .b(weight_2_11_reg[1]), .cin(weight_2_11_reg[2]), .sum(weight_3_11[1]), .cout(weight_3_12[0]));
full_adder fa518(.a(weight_2_12_reg[0]), .b(weight_2_12_reg[1]), .cin(weight_2_12_reg[2]), .sum(weight_3_12[1]), .cout(weight_3_13[0]));
full_adder fa519(.a(weight_2_13_reg[0]), .b(weight_2_13_reg[1]), .cin(weight_2_13_reg[2]), .sum(weight_3_13[1]), .cout(weight_3_14[0]));
full_adder fa520(.a(weight_2_14_reg[0]), .b(weight_2_14_reg[1]), .cin(weight_2_14_reg[2]), .sum(weight_3_14[1]), .cout(weight_3_15[0]));
full_adder fa521(.a(weight_2_15_reg[0]), .b(weight_2_15_reg[1]), .cin(weight_2_15_reg[2]), .sum(weight_3_15[1]), .cout(weight_3_16[0]));
full_adder fa522(.a(weight_2_16_reg[0]), .b(weight_2_16_reg[1]), .cin(weight_2_16_reg[2]), .sum(weight_3_16[1]), .cout(weight_3_17[0]));
full_adder fa523(.a(weight_2_17_reg[0]), .b(weight_2_17_reg[1]), .cin(weight_2_17_reg[2]), .sum(weight_3_17[1]), .cout(weight_3_18[0]));
full_adder fa524(.a(weight_2_18_reg[0]), .b(weight_2_18_reg[1]), .cin(weight_2_18_reg[2]), .sum(weight_3_18[1]), .cout(weight_3_19[0]));
full_adder fa525(.a(weight_2_19_reg[0]), .b(weight_2_19_reg[1]), .cin(weight_2_19_reg[2]), .sum(weight_3_19[1]), .cout(weight_3_20[0]));
full_adder fa526(.a(weight_2_20_reg[0]), .b(weight_2_20_reg[1]), .cin(weight_2_20_reg[2]), .sum(weight_3_20[1]), .cout(weight_3_21[0]));
full_adder fa527(.a(weight_2_21_reg[0]), .b(weight_2_21_reg[1]), .cin(weight_2_21_reg[2]), .sum(weight_3_21[1]), .cout(weight_3_22[0]));
full_adder fa528(.a(weight_2_22_reg[0]), .b(weight_2_22_reg[1]), .cin(weight_2_22_reg[2]), .sum(weight_3_22[1]), .cout(weight_3_23[0]));
full_adder fa529(.a(weight_2_23_reg[0]), .b(weight_2_23_reg[1]), .cin(weight_2_23_reg[2]), .sum(weight_3_23[1]), .cout(weight_3_24[0]));
full_adder fa530(.a(weight_2_24_reg[0]), .b(weight_2_24_reg[1]), .cin(weight_2_24_reg[2]), .sum(weight_3_24[1]), .cout(weight_3_25[0]));
full_adder fa531(.a(weight_2_25_reg[0]), .b(weight_2_25_reg[1]), .cin(weight_2_25_reg[2]), .sum(weight_3_25[1]), .cout(weight_3_26[0]));
full_adder fa532(.a(weight_2_26_reg[0]), .b(weight_2_26_reg[1]), .cin(weight_2_26_reg[2]), .sum(weight_3_26[1]), .cout(weight_3_27[0]));
full_adder fa533(.a(weight_2_27_reg[0]), .b(weight_2_27_reg[1]), .cin(weight_2_27_reg[2]), .sum(weight_3_27[1]), .cout(weight_3_28[0]));
full_adder fa534(.a(weight_2_28_reg[0]), .b(weight_2_28_reg[1]), .cin(weight_2_28_reg[2]), .sum(weight_3_28[1]), .cout(weight_3_29[0]));
full_adder fa535(.a(weight_2_29_reg[0]), .b(weight_2_29_reg[1]), .cin(weight_2_29_reg[2]), .sum(weight_3_29[1]), .cout(weight_3_30[0]));
full_adder fa536(.a(weight_2_30_reg[0]), .b(weight_2_30_reg[1]), .cin(weight_2_30_reg[2]), .sum(weight_3_30[1]), .cout(weight_3_31[0]));
full_adder fa537(.a(weight_2_31_reg[0]), .b(weight_2_31_reg[1]), .cin(weight_2_31_reg[2]), .sum(weight_3_31[1]), .cout(weight_3_32[0]));
full_adder fa538(.a(weight_2_32_reg[0]), .b(weight_2_32_reg[1]), .cin(weight_2_32_reg[2]), .sum(weight_3_32[1]), .cout(weight_3_33[0]));
full_adder fa539(.a(weight_2_33_reg[0]), .b(weight_2_33_reg[1]), .cin(weight_2_33_reg[2]), .sum(weight_3_33[1]), .cout(weight_3_34[0]));
full_adder fa540(.a(weight_2_34_reg[0]), .b(weight_2_34_reg[1]), .cin(weight_2_34_reg[2]), .sum(weight_3_34[1]), .cout(weight_3_35[0]));
half_adder ha41(.a(weight_2_35_reg[0]), .b(weight_2_35_reg[1]), .sum(weight_3_35[1]), .cout(weight_3_36[0]));
half_adder ha42(.a(weight_2_36_reg[0]), .b(weight_2_36_reg[1]), .sum(weight_3_36[1]), .cout(weight_3_37[0]));
assign weight_3_37[1] = weight_2_37_reg[0];
assign weight_3_38[0] = weight_2_38_reg[0];
assign weight_3_39[0] = weight_2_39_reg[0];
assign weight_3_7[2] = weight_2_7_reg[3];
assign weight_3_8[2] = weight_2_8_reg[3];
half_adder ha43(.a(weight_2_9_reg[3]), .b(weight_2_9_reg[4]), .sum(weight_3_9[2]), .cout(weight_3_10[2]));
half_adder ha44(.a(weight_2_10_reg[3]), .b(weight_2_10_reg[4]), .sum(weight_3_10[3]), .cout(weight_3_11[2]));
half_adder ha45(.a(weight_2_11_reg[3]), .b(weight_2_11_reg[4]), .sum(weight_3_11[3]), .cout(weight_3_12[2]));
full_adder fa541(.a(weight_2_12_reg[3]), .b(weight_2_12_reg[4]), .cin(weight_2_12_reg[5]), .sum(weight_3_12[3]), .cout(weight_3_13[2]));
full_adder fa542(.a(weight_2_13_reg[3]), .b(weight_2_13_reg[4]), .cin(weight_2_13_reg[5]), .sum(weight_3_13[3]), .cout(weight_3_14[2]));
full_adder fa543(.a(weight_2_14_reg[3]), .b(weight_2_14_reg[4]), .cin(weight_2_14_reg[5]), .sum(weight_3_14[3]), .cout(weight_3_15[2]));
full_adder fa544(.a(weight_2_15_reg[3]), .b(weight_2_15_reg[4]), .cin(weight_2_15_reg[5]), .sum(weight_3_15[3]), .cout(weight_3_16[2]));
full_adder fa545(.a(weight_2_16_reg[3]), .b(weight_2_16_reg[4]), .cin(weight_2_16_reg[5]), .sum(weight_3_16[3]), .cout(weight_3_17[2]));
full_adder fa546(.a(weight_2_17_reg[3]), .b(weight_2_17_reg[4]), .cin(weight_2_17_reg[5]), .sum(weight_3_17[3]), .cout(weight_3_18[2]));
full_adder fa547(.a(weight_2_18_reg[3]), .b(weight_2_18_reg[4]), .cin(weight_2_18_reg[5]), .sum(weight_3_18[3]), .cout(weight_3_19[2]));
full_adder fa548(.a(weight_2_19_reg[3]), .b(weight_2_19_reg[4]), .cin(weight_2_19_reg[5]), .sum(weight_3_19[3]), .cout(weight_3_20[2]));
full_adder fa549(.a(weight_2_20_reg[3]), .b(weight_2_20_reg[4]), .cin(weight_2_20_reg[5]), .sum(weight_3_20[3]), .cout(weight_3_21[2]));
full_adder fa550(.a(weight_2_21_reg[3]), .b(weight_2_21_reg[4]), .cin(weight_2_21_reg[5]), .sum(weight_3_21[3]), .cout(weight_3_22[2]));
full_adder fa551(.a(weight_2_22_reg[3]), .b(weight_2_22_reg[4]), .cin(weight_2_22_reg[5]), .sum(weight_3_22[3]), .cout(weight_3_23[2]));
full_adder fa552(.a(weight_2_23_reg[3]), .b(weight_2_23_reg[4]), .cin(weight_2_23_reg[5]), .sum(weight_3_23[3]), .cout(weight_3_24[2]));
full_adder fa553(.a(weight_2_24_reg[3]), .b(weight_2_24_reg[4]), .cin(weight_2_24_reg[5]), .sum(weight_3_24[3]), .cout(weight_3_25[2]));
full_adder fa554(.a(weight_2_25_reg[3]), .b(weight_2_25_reg[4]), .cin(weight_2_25_reg[5]), .sum(weight_3_25[3]), .cout(weight_3_26[2]));
full_adder fa555(.a(weight_2_26_reg[3]), .b(weight_2_26_reg[4]), .cin(weight_2_26_reg[5]), .sum(weight_3_26[3]), .cout(weight_3_27[2]));
full_adder fa556(.a(weight_2_27_reg[3]), .b(weight_2_27_reg[4]), .cin(weight_2_27_reg[5]), .sum(weight_3_27[3]), .cout(weight_3_28[2]));
full_adder fa557(.a(weight_2_28_reg[3]), .b(weight_2_28_reg[4]), .cin(weight_2_28_reg[5]), .sum(weight_3_28[3]), .cout(weight_3_29[2]));
full_adder fa558(.a(weight_2_29_reg[3]), .b(weight_2_29_reg[4]), .cin(weight_2_29_reg[5]), .sum(weight_3_29[3]), .cout(weight_3_30[2]));
full_adder fa559(.a(weight_2_30_reg[3]), .b(weight_2_30_reg[4]), .cin(weight_2_30_reg[5]), .sum(weight_3_30[3]), .cout(weight_3_31[2]));
full_adder fa560(.a(weight_2_31_reg[3]), .b(weight_2_31_reg[4]), .cin(weight_2_31_reg[5]), .sum(weight_3_31[3]), .cout(weight_3_32[2]));
full_adder fa561(.a(weight_2_32_reg[3]), .b(weight_2_32_reg[4]), .cin(weight_2_32_reg[5]), .sum(weight_3_32[3]), .cout(weight_3_33[2]));
full_adder fa562(.a(weight_2_33_reg[3]), .b(weight_2_33_reg[4]), .cin(weight_2_33_reg[5]), .sum(weight_3_33[3]), .cout(weight_3_34[2]));
full_adder fa563(.a(weight_2_34_reg[3]), .b(weight_2_34_reg[4]), .cin(weight_2_34_reg[5]), .sum(weight_3_34[3]), .cout(weight_3_35[2]));
full_adder fa564(.a(weight_2_35_reg[2]), .b(weight_2_35_reg[3]), .cin(weight_2_35_reg[4]), .sum(weight_3_35[3]), .cout(weight_3_36[2]));
full_adder fa565(.a(weight_2_36_reg[2]), .b(weight_2_36_reg[3]), .cin(weight_2_36_reg[4]), .sum(weight_3_36[3]), .cout(weight_3_37[2]));
full_adder fa566(.a(weight_2_37_reg[1]), .b(weight_2_37_reg[2]), .cin(weight_2_37_reg[3]), .sum(weight_3_37[3]), .cout(weight_3_38[1]));
full_adder fa567(.a(weight_2_38_reg[1]), .b(weight_2_38_reg[2]), .cin(weight_2_38_reg[3]), .sum(weight_3_38[2]), .cout(weight_3_39[1]));
full_adder fa568(.a(weight_2_39_reg[1]), .b(weight_2_39_reg[2]), .cin(weight_2_39_reg[3]), .sum(weight_3_39[2]), .cout(weight_3_40[0]));
full_adder fa569(.a(weight_2_40_reg[0]), .b(weight_2_40_reg[1]), .cin(weight_2_40_reg[2]), .sum(weight_3_40[1]), .cout(weight_3_41[0]));
half_adder ha46(.a(weight_2_41_reg[0]), .b(weight_2_41_reg[1]), .sum(weight_3_41[1]), .cout(weight_3_42[0]));
half_adder ha47(.a(weight_2_42_reg[0]), .b(weight_2_42_reg[1]), .sum(weight_3_42[1]), .cout(weight_3_43[0]));
half_adder ha48(.a(weight_2_43_reg[0]), .b(weight_2_43_reg[1]), .sum(weight_3_43[1]), .cout(weight_3_44[0]));
assign weight_3_44[1] = weight_2_44_reg[0];
assign weight_3_45[0] = weight_2_45_reg[0];
assign weight_3_14[4] = weight_2_14_reg[6];
assign weight_3_15[4] = weight_2_15_reg[6];
half_adder ha49(.a(weight_2_16_reg[6]), .b(weight_2_16_reg[7]), .sum(weight_3_16[4]), .cout(weight_3_17[4]));
half_adder ha50(.a(weight_2_17_reg[6]), .b(weight_2_17_reg[7]), .sum(weight_3_17[5]), .cout(weight_3_18[4]));
full_adder fa570(.a(weight_2_18_reg[6]), .b(weight_2_18_reg[7]), .cin(weight_2_18_reg[8]), .sum(weight_3_18[5]), .cout(weight_3_19[4]));
full_adder fa571(.a(weight_2_19_reg[6]), .b(weight_2_19_reg[7]), .cin(weight_2_19_reg[8]), .sum(weight_3_19[5]), .cout(weight_3_20[4]));
full_adder fa572(.a(weight_2_20_reg[6]), .b(weight_2_20_reg[7]), .cin(weight_2_20_reg[8]), .sum(weight_3_20[5]), .cout(weight_3_21[4]));
full_adder fa573(.a(weight_2_21_reg[6]), .b(weight_2_21_reg[7]), .cin(weight_2_21_reg[8]), .sum(weight_3_21[5]), .cout(weight_3_22[4]));
full_adder fa574(.a(weight_2_22_reg[6]), .b(weight_2_22_reg[7]), .cin(weight_2_22_reg[8]), .sum(weight_3_22[5]), .cout(weight_3_23[4]));
full_adder fa575(.a(weight_2_23_reg[6]), .b(weight_2_23_reg[7]), .cin(weight_2_23_reg[8]), .sum(weight_3_23[5]), .cout(weight_3_24[4]));
full_adder fa576(.a(weight_2_24_reg[6]), .b(weight_2_24_reg[7]), .cin(weight_2_24_reg[8]), .sum(weight_3_24[5]), .cout(weight_3_25[4]));
full_adder fa577(.a(weight_2_25_reg[6]), .b(weight_2_25_reg[7]), .cin(weight_2_25_reg[8]), .sum(weight_3_25[5]), .cout(weight_3_26[4]));
full_adder fa578(.a(weight_2_26_reg[6]), .b(weight_2_26_reg[7]), .cin(weight_2_26_reg[8]), .sum(weight_3_26[5]), .cout(weight_3_27[4]));
full_adder fa579(.a(weight_2_27_reg[6]), .b(weight_2_27_reg[7]), .cin(weight_2_27_reg[8]), .sum(weight_3_27[5]), .cout(weight_3_28[4]));
full_adder fa580(.a(weight_2_28_reg[6]), .b(weight_2_28_reg[7]), .cin(weight_2_28_reg[8]), .sum(weight_3_28[5]), .cout(weight_3_29[4]));
full_adder fa581(.a(weight_2_29_reg[6]), .b(weight_2_29_reg[7]), .cin(weight_2_29_reg[8]), .sum(weight_3_29[5]), .cout(weight_3_30[4]));
full_adder fa582(.a(weight_2_30_reg[6]), .b(weight_2_30_reg[7]), .cin(weight_2_30_reg[8]), .sum(weight_3_30[5]), .cout(weight_3_31[4]));
full_adder fa583(.a(weight_2_31_reg[6]), .b(weight_2_31_reg[7]), .cin(weight_2_31_reg[8]), .sum(weight_3_31[5]), .cout(weight_3_32[4]));
full_adder fa584(.a(weight_2_32_reg[6]), .b(weight_2_32_reg[7]), .cin(weight_2_32_reg[8]), .sum(weight_3_32[5]), .cout(weight_3_33[4]));
full_adder fa585(.a(weight_2_33_reg[6]), .b(weight_2_33_reg[7]), .cin(weight_2_33_reg[8]), .sum(weight_3_33[5]), .cout(weight_3_34[4]));
full_adder fa586(.a(weight_2_34_reg[6]), .b(weight_2_34_reg[7]), .cin(weight_2_34_reg[8]), .sum(weight_3_34[5]), .cout(weight_3_35[4]));
full_adder fa587(.a(weight_2_35_reg[5]), .b(weight_2_35_reg[6]), .cin(weight_2_35_reg[7]), .sum(weight_3_35[5]), .cout(weight_3_36[4]));
full_adder fa588(.a(weight_2_36_reg[5]), .b(weight_2_36_reg[6]), .cin(weight_2_36_reg[7]), .sum(weight_3_36[5]), .cout(weight_3_37[4]));
full_adder fa589(.a(weight_2_37_reg[4]), .b(weight_2_37_reg[5]), .cin(weight_2_37_reg[6]), .sum(weight_3_37[5]), .cout(weight_3_38[3]));
full_adder fa590(.a(weight_2_38_reg[4]), .b(weight_2_38_reg[5]), .cin(weight_2_38_reg[6]), .sum(weight_3_38[4]), .cout(weight_3_39[3]));
full_adder fa591(.a(weight_2_39_reg[4]), .b(weight_2_39_reg[5]), .cin(weight_2_39_reg[6]), .sum(weight_3_39[4]), .cout(weight_3_40[2]));
full_adder fa592(.a(weight_2_40_reg[3]), .b(weight_2_40_reg[4]), .cin(weight_2_40_reg[5]), .sum(weight_3_40[3]), .cout(weight_3_41[2]));
full_adder fa593(.a(weight_2_41_reg[2]), .b(weight_2_41_reg[3]), .cin(weight_2_41_reg[4]), .sum(weight_3_41[3]), .cout(weight_3_42[2]));
full_adder fa594(.a(weight_2_42_reg[2]), .b(weight_2_42_reg[3]), .cin(weight_2_42_reg[4]), .sum(weight_3_42[3]), .cout(weight_3_43[2]));
full_adder fa595(.a(weight_2_43_reg[2]), .b(weight_2_43_reg[3]), .cin(weight_2_43_reg[4]), .sum(weight_3_43[3]), .cout(weight_3_44[2]));
full_adder fa596(.a(weight_2_44_reg[1]), .b(weight_2_44_reg[2]), .cin(weight_2_44_reg[3]), .sum(weight_3_44[3]), .cout(weight_3_45[1]));
full_adder fa597(.a(weight_2_45_reg[1]), .b(weight_2_45_reg[2]), .cin(weight_2_45_reg[3]), .sum(weight_3_45[2]), .cout(weight_3_46[0]));
full_adder fa598(.a(weight_2_46_reg[0]), .b(weight_2_46_reg[1]), .cin(weight_2_46_reg[2]), .sum(weight_3_46[1]), .cout(weight_3_47[0]));
full_adder fa599(.a(weight_2_47_reg[0]), .b(weight_2_47_reg[1]), .cin(weight_2_47_reg[2]), .sum(weight_3_47[1]), .cout(weight_3_48[0]));
full_adder fa600(.a(weight_2_48_reg[0]), .b(weight_2_48_reg[1]), .cin(weight_2_48_reg[2]), .sum(weight_3_48[1]), .cout(weight_3_49[0]));
half_adder ha51(.a(weight_2_49_reg[0]), .b(weight_2_49_reg[1]), .sum(weight_3_49[1]), .cout(weight_3_50[0]));
assign weight_3_50[1] = weight_2_50_reg[0];
assign weight_3_51[0] = weight_2_51_reg[0];
assign weight_3_52[0] = weight_2_52_reg[0];
assign weight_3_21[6] = weight_2_21_reg[9];
assign weight_3_22[6] = weight_2_22_reg[9];
half_adder ha52(.a(weight_2_23_reg[9]), .b(weight_2_23_reg[10]), .sum(weight_3_23[6]), .cout(weight_3_24[6]));
half_adder ha53(.a(weight_2_24_reg[9]), .b(weight_2_24_reg[10]), .sum(weight_3_24[7]), .cout(weight_3_25[6]));
full_adder fa601(.a(weight_2_25_reg[9]), .b(weight_2_25_reg[10]), .cin(weight_2_25_reg[11]), .sum(weight_3_25[7]), .cout(weight_3_26[6]));
full_adder fa602(.a(weight_2_26_reg[9]), .b(weight_2_26_reg[10]), .cin(weight_2_26_reg[11]), .sum(weight_3_26[7]), .cout(weight_3_27[6]));
full_adder fa603(.a(weight_2_27_reg[9]), .b(weight_2_27_reg[10]), .cin(weight_2_27_reg[11]), .sum(weight_3_27[7]), .cout(weight_3_28[6]));
full_adder fa604(.a(weight_2_28_reg[9]), .b(weight_2_28_reg[10]), .cin(weight_2_28_reg[11]), .sum(weight_3_28[7]), .cout(weight_3_29[6]));
full_adder fa605(.a(weight_2_29_reg[9]), .b(weight_2_29_reg[10]), .cin(weight_2_29_reg[11]), .sum(weight_3_29[7]), .cout(weight_3_30[6]));
full_adder fa606(.a(weight_2_30_reg[9]), .b(weight_2_30_reg[10]), .cin(weight_2_30_reg[11]), .sum(weight_3_30[7]), .cout(weight_3_31[6]));
full_adder fa607(.a(weight_2_31_reg[9]), .b(weight_2_31_reg[10]), .cin(weight_2_31_reg[11]), .sum(weight_3_31[7]), .cout(weight_3_32[6]));
full_adder fa608(.a(weight_2_32_reg[9]), .b(weight_2_32_reg[10]), .cin(weight_2_32_reg[11]), .sum(weight_3_32[7]), .cout(weight_3_33[6]));
full_adder fa609(.a(weight_2_33_reg[9]), .b(weight_2_33_reg[10]), .cin(weight_2_33_reg[11]), .sum(weight_3_33[7]), .cout(weight_3_34[6]));
full_adder fa610(.a(weight_2_34_reg[9]), .b(weight_2_34_reg[10]), .cin(weight_2_34_reg[11]), .sum(weight_3_34[7]), .cout(weight_3_35[6]));
full_adder fa611(.a(weight_2_35_reg[8]), .b(weight_2_35_reg[9]), .cin(weight_2_35_reg[10]), .sum(weight_3_35[7]), .cout(weight_3_36[6]));
full_adder fa612(.a(weight_2_36_reg[8]), .b(weight_2_36_reg[9]), .cin(weight_2_36_reg[10]), .sum(weight_3_36[7]), .cout(weight_3_37[6]));
full_adder fa613(.a(weight_2_37_reg[7]), .b(weight_2_37_reg[8]), .cin(weight_2_37_reg[9]), .sum(weight_3_37[7]), .cout(weight_3_38[5]));
full_adder fa614(.a(weight_2_38_reg[7]), .b(weight_2_38_reg[8]), .cin(weight_2_38_reg[9]), .sum(weight_3_38[6]), .cout(weight_3_39[5]));
full_adder fa615(.a(weight_2_39_reg[7]), .b(weight_2_39_reg[8]), .cin(weight_2_39_reg[9]), .sum(weight_3_39[6]), .cout(weight_3_40[4]));
full_adder fa616(.a(weight_2_40_reg[6]), .b(weight_2_40_reg[7]), .cin(weight_2_40_reg[8]), .sum(weight_3_40[5]), .cout(weight_3_41[4]));
full_adder fa617(.a(weight_2_41_reg[5]), .b(weight_2_41_reg[6]), .cin(weight_2_41_reg[7]), .sum(weight_3_41[5]), .cout(weight_3_42[4]));
full_adder fa618(.a(weight_2_42_reg[5]), .b(weight_2_42_reg[6]), .cin(weight_2_42_reg[7]), .sum(weight_3_42[5]), .cout(weight_3_43[4]));
full_adder fa619(.a(weight_2_43_reg[5]), .b(weight_2_43_reg[6]), .cin(weight_2_43_reg[7]), .sum(weight_3_43[5]), .cout(weight_3_44[4]));
full_adder fa620(.a(weight_2_44_reg[4]), .b(weight_2_44_reg[5]), .cin(weight_2_44_reg[6]), .sum(weight_3_44[5]), .cout(weight_3_45[3]));
full_adder fa621(.a(weight_2_45_reg[4]), .b(weight_2_45_reg[5]), .cin(weight_2_45_reg[6]), .sum(weight_3_45[4]), .cout(weight_3_46[2]));
full_adder fa622(.a(weight_2_46_reg[3]), .b(weight_2_46_reg[4]), .cin(weight_2_46_reg[5]), .sum(weight_3_46[3]), .cout(weight_3_47[2]));
full_adder fa623(.a(weight_2_47_reg[3]), .b(weight_2_47_reg[4]), .cin(weight_2_47_reg[5]), .sum(weight_3_47[3]), .cout(weight_3_48[2]));
full_adder fa624(.a(weight_2_48_reg[3]), .b(weight_2_48_reg[4]), .cin(weight_2_48_reg[5]), .sum(weight_3_48[3]), .cout(weight_3_49[2]));
full_adder fa625(.a(weight_2_49_reg[2]), .b(weight_2_49_reg[3]), .cin(weight_2_49_reg[4]), .sum(weight_3_49[3]), .cout(weight_3_50[2]));
full_adder fa626(.a(weight_2_50_reg[1]), .b(weight_2_50_reg[2]), .cin(weight_2_50_reg[3]), .sum(weight_3_50[3]), .cout(weight_3_51[1]));
full_adder fa627(.a(weight_2_51_reg[1]), .b(weight_2_51_reg[2]), .cin(weight_2_51_reg[3]), .sum(weight_3_51[2]), .cout(weight_3_52[1]));
full_adder fa628(.a(weight_2_52_reg[1]), .b(weight_2_52_reg[2]), .cin(weight_2_52_reg[3]), .sum(weight_3_52[2]), .cout(weight_3_53[0]));
full_adder fa629(.a(weight_2_53_reg[0]), .b(weight_2_53_reg[1]), .cin(weight_2_53_reg[2]), .sum(weight_3_53[1]), .cout(weight_3_54[0]));
full_adder fa630(.a(weight_2_54_reg[0]), .b(weight_2_54_reg[1]), .cin(weight_2_54_reg[2]), .sum(weight_3_54[1]), .cout(weight_3_55[0]));
half_adder ha54(.a(weight_2_55_reg[0]), .b(weight_2_55_reg[1]), .sum(weight_3_55[1]), .cout(weight_3_56[0]));
half_adder ha55(.a(weight_2_56_reg[0]), .b(weight_2_56_reg[1]), .sum(weight_3_56[1]), .cout(weight_3_57[0]));
half_adder ha56(.a(weight_2_57_reg[0]), .b(weight_2_57_reg[1]), .sum(weight_3_57[1]), .cout(weight_3_58[0]));
assign weight_3_58[1] = weight_2_58_reg[0];
assign weight_3_27[8] = weight_2_27_reg[12];
assign weight_3_28[8] = weight_2_28_reg[12];
assign weight_3_29[8] = weight_2_29_reg[12];
half_adder ha57(.a(weight_2_30_reg[12]), .b(weight_2_30_reg[13]), .sum(weight_3_30[8]), .cout(weight_3_31[8]));
full_adder fa631(.a(weight_2_31_reg[12]), .b(weight_2_31_reg[13]), .cin(weight_2_31_reg[14]), .sum(weight_3_31[9]), .cout(weight_3_32[8]));
full_adder fa632(.a(weight_2_32_reg[12]), .b(weight_2_32_reg[13]), .cin(weight_2_32_reg[14]), .sum(weight_3_32[9]), .cout(weight_3_33[8]));
full_adder fa633(.a(weight_2_33_reg[12]), .b(weight_2_33_reg[13]), .cin(weight_2_33_reg[14]), .sum(weight_3_33[9]), .cout(weight_3_34[8]));
full_adder fa634(.a(weight_2_34_reg[12]), .b(weight_2_34_reg[13]), .cin(weight_2_34_reg[14]), .sum(weight_3_34[9]), .cout(weight_3_35[8]));
full_adder fa635(.a(weight_2_35_reg[11]), .b(weight_2_35_reg[12]), .cin(weight_2_35_reg[13]), .sum(weight_3_35[9]), .cout(weight_3_36[8]));
full_adder fa636(.a(weight_2_36_reg[11]), .b(weight_2_36_reg[12]), .cin(weight_2_36_reg[13]), .sum(weight_3_36[9]), .cout(weight_3_37[8]));
full_adder fa637(.a(weight_2_37_reg[10]), .b(weight_2_37_reg[11]), .cin(weight_2_37_reg[12]), .sum(weight_3_37[9]), .cout(weight_3_38[7]));
full_adder fa638(.a(weight_2_38_reg[10]), .b(weight_2_38_reg[11]), .cin(weight_2_38_reg[12]), .sum(weight_3_38[8]), .cout(weight_3_39[7]));
full_adder fa639(.a(weight_2_39_reg[10]), .b(weight_2_39_reg[11]), .cin(weight_2_39_reg[12]), .sum(weight_3_39[8]), .cout(weight_3_40[6]));
full_adder fa640(.a(weight_2_40_reg[9]), .b(weight_2_40_reg[10]), .cin(weight_2_40_reg[11]), .sum(weight_3_40[7]), .cout(weight_3_41[6]));
full_adder fa641(.a(weight_2_41_reg[8]), .b(weight_2_41_reg[9]), .cin(weight_2_41_reg[10]), .sum(weight_3_41[7]), .cout(weight_3_42[6]));
full_adder fa642(.a(weight_2_42_reg[8]), .b(weight_2_42_reg[9]), .cin(weight_2_42_reg[10]), .sum(weight_3_42[7]), .cout(weight_3_43[6]));
full_adder fa643(.a(weight_2_43_reg[8]), .b(weight_2_43_reg[9]), .cin(weight_2_43_reg[10]), .sum(weight_3_43[7]), .cout(weight_3_44[6]));
full_adder fa644(.a(weight_2_44_reg[7]), .b(weight_2_44_reg[8]), .cin(weight_2_44_reg[9]), .sum(weight_3_44[7]), .cout(weight_3_45[5]));
full_adder fa645(.a(weight_2_45_reg[7]), .b(weight_2_45_reg[8]), .cin(weight_2_45_reg[9]), .sum(weight_3_45[6]), .cout(weight_3_46[4]));
full_adder fa646(.a(weight_2_46_reg[6]), .b(weight_2_46_reg[7]), .cin(weight_2_46_reg[8]), .sum(weight_3_46[5]), .cout(weight_3_47[4]));
full_adder fa647(.a(weight_2_47_reg[6]), .b(weight_2_47_reg[7]), .cin(weight_2_47_reg[8]), .sum(weight_3_47[5]), .cout(weight_3_48[4]));
full_adder fa648(.a(weight_2_48_reg[6]), .b(weight_2_48_reg[7]), .cin(weight_2_48_reg[8]), .sum(weight_3_48[5]), .cout(weight_3_49[4]));
full_adder fa649(.a(weight_2_49_reg[5]), .b(weight_2_49_reg[6]), .cin(weight_2_49_reg[7]), .sum(weight_3_49[5]), .cout(weight_3_50[4]));
full_adder fa650(.a(weight_2_50_reg[4]), .b(weight_2_50_reg[5]), .cin(weight_2_50_reg[6]), .sum(weight_3_50[5]), .cout(weight_3_51[3]));
full_adder fa651(.a(weight_2_51_reg[4]), .b(weight_2_51_reg[5]), .cin(weight_2_51_reg[6]), .sum(weight_3_51[4]), .cout(weight_3_52[3]));
full_adder fa652(.a(weight_2_52_reg[4]), .b(weight_2_52_reg[5]), .cin(weight_2_52_reg[6]), .sum(weight_3_52[4]), .cout(weight_3_53[2]));
full_adder fa653(.a(weight_2_53_reg[3]), .b(weight_2_53_reg[4]), .cin(weight_2_53_reg[5]), .sum(weight_3_53[3]), .cout(weight_3_54[2]));
full_adder fa654(.a(weight_2_54_reg[3]), .b(weight_2_54_reg[4]), .cin(weight_2_54_reg[5]), .sum(weight_3_54[3]), .cout(weight_3_55[2]));
full_adder fa655(.a(weight_2_55_reg[2]), .b(weight_2_55_reg[3]), .cin(weight_2_55_reg[4]), .sum(weight_3_55[3]), .cout(weight_3_56[2]));
full_adder fa656(.a(weight_2_56_reg[2]), .b(weight_2_56_reg[3]), .cin(weight_2_56_reg[4]), .sum(weight_3_56[3]), .cout(weight_3_57[2]));
full_adder fa657(.a(weight_2_57_reg[2]), .b(weight_2_57_reg[3]), .cin(weight_2_57_reg[4]), .sum(weight_3_57[3]), .cout(weight_3_58[2]));
full_adder fa658(.a(weight_2_58_reg[1]), .b(weight_2_58_reg[2]), .cin(weight_2_58_reg[3]), .sum(weight_3_58[3]), .cout(weight_3_59[0]));
full_adder fa659(.a(weight_2_59_reg[0]), .b(weight_2_59_reg[1]), .cin(weight_2_59_reg[2]), .sum(weight_3_59[1]), .cout(weight_3_60[0]));
full_adder fa660(.a(weight_2_60_reg[0]), .b(weight_2_60_reg[1]), .cin(weight_2_60_reg[2]), .sum(weight_3_60[1]), .cout(weight_3_61[0]));
full_adder fa661(.a(weight_2_61_reg[0]), .b(weight_2_61_reg[1]), .cin(weight_2_61_reg[2]), .sum(weight_3_61[1]), .cout(weight_3_62[0]));
assign weight_3_62[1] = weight_2_62_reg;
logic weight_4_0;
logic weight_4_1;
logic weight_4_2;
logic weight_4_3;
logic weight_4_4;
logic [1:0] weight_4_5;
logic [1:0] weight_4_6;
logic [1:0] weight_4_7;
logic [1:0] weight_4_8;
logic [1:0] weight_4_9;
logic [2:0] weight_4_10;
logic [2:0] weight_4_11;
logic [2:0] weight_4_12;
logic [2:0] weight_4_13;
logic [2:0] weight_4_14;
logic [3:0] weight_4_15;
logic [3:0] weight_4_16;
logic [3:0] weight_4_17;
logic [3:0] weight_4_18;
logic [3:0] weight_4_19;
logic [3:0] weight_4_20;
logic [4:0] weight_4_21;
logic [4:0] weight_4_22;
logic [4:0] weight_4_23;
logic [4:0] weight_4_24;
logic [5:0] weight_4_25;
logic [5:0] weight_4_26;
logic [5:0] weight_4_27;
logic [5:0] weight_4_28;
logic [5:0] weight_4_29;
logic [5:0] weight_4_30;
logic [6:0] weight_4_31;
logic [6:0] weight_4_32;
logic [6:0] weight_4_33;
logic [6:0] weight_4_34;
logic [6:0] weight_4_35;
logic [6:0] weight_4_36;
logic [6:0] weight_4_37;
logic [6:0] weight_4_38;
logic [6:0] weight_4_39;
logic [6:0] weight_4_40;
logic [5:0] weight_4_41;
logic [5:0] weight_4_42;
logic [5:0] weight_4_43;
logic [5:0] weight_4_44;
logic [4:0] weight_4_45;
logic [4:0] weight_4_46;
logic [4:0] weight_4_47;
logic [4:0] weight_4_48;
logic [4:0] weight_4_49;
logic [4:0] weight_4_50;
logic [4:0] weight_4_51;
logic [3:0] weight_4_52;
logic [2:0] weight_4_53;
logic [2:0] weight_4_54;
logic [2:0] weight_4_55;
logic [2:0] weight_4_56;
logic [2:0] weight_4_57;
logic [2:0] weight_4_58;
logic [2:0] weight_4_59;
logic [1:0] weight_4_60;
logic [1:0] weight_4_61;
logic [1:0] weight_4_62;

logic en_reg_2;
logic weight_4_0_reg;
logic weight_4_1_reg;
logic weight_4_2_reg;
logic weight_4_3_reg;
logic weight_4_4_reg;
logic [1:0] weight_4_5_reg;
logic [1:0] weight_4_6_reg;
logic [1:0] weight_4_7_reg;
logic [1:0] weight_4_8_reg;
logic [1:0] weight_4_9_reg;
logic [2:0] weight_4_10_reg;
logic [2:0] weight_4_11_reg;
logic [2:0] weight_4_12_reg;
logic [2:0] weight_4_13_reg;
logic [2:0] weight_4_14_reg;
logic [3:0] weight_4_15_reg;
logic [3:0] weight_4_16_reg;
logic [3:0] weight_4_17_reg;
logic [3:0] weight_4_18_reg;
logic [3:0] weight_4_19_reg;
logic [3:0] weight_4_20_reg;
logic [4:0] weight_4_21_reg;
logic [4:0] weight_4_22_reg;
logic [4:0] weight_4_23_reg;
logic [4:0] weight_4_24_reg;
logic [5:0] weight_4_25_reg;
logic [5:0] weight_4_26_reg;
logic [5:0] weight_4_27_reg;
logic [5:0] weight_4_28_reg;
logic [5:0] weight_4_29_reg;
logic [5:0] weight_4_30_reg;
logic [6:0] weight_4_31_reg;
logic [6:0] weight_4_32_reg;
logic [6:0] weight_4_33_reg;
logic [6:0] weight_4_34_reg;
logic [6:0] weight_4_35_reg;
logic [6:0] weight_4_36_reg;
logic [6:0] weight_4_37_reg;
logic [6:0] weight_4_38_reg;
logic [6:0] weight_4_39_reg;
logic [6:0] weight_4_40_reg;
logic [5:0] weight_4_41_reg;
logic [5:0] weight_4_42_reg;
logic [5:0] weight_4_43_reg;
logic [5:0] weight_4_44_reg;
logic [4:0] weight_4_45_reg;
logic [4:0] weight_4_46_reg;
logic [4:0] weight_4_47_reg;
logic [4:0] weight_4_48_reg;
logic [4:0] weight_4_49_reg;
logic [4:0] weight_4_50_reg;
logic [4:0] weight_4_51_reg;
logic [3:0] weight_4_52_reg;
logic [2:0] weight_4_53_reg;
logic [2:0] weight_4_54_reg;
logic [2:0] weight_4_55_reg;
logic [2:0] weight_4_56_reg;
logic [2:0] weight_4_57_reg;
logic [2:0] weight_4_58_reg;
logic [2:0] weight_4_59_reg;
logic [1:0] weight_4_60_reg;
logic [1:0] weight_4_61_reg;
logic [1:0] weight_4_62_reg;

// Second pipeline stage
always_ff @(posedge clk, negedge nrst) begin
    if (~nrst | multiplier_if.ready) begin
        en_reg_2 <= '0;
        weight_4_0_reg <= '0;
        weight_4_1_reg <= '0;
        weight_4_2_reg <= '0;
        weight_4_3_reg <= '0;
        weight_4_4_reg <= '0;
        weight_4_5_reg <= '0;
        weight_4_6_reg <= '0;
        weight_4_7_reg <= '0;
        weight_4_8_reg <= '0;
        weight_4_9_reg <= '0;
        weight_4_10_reg <= '0;
        weight_4_11_reg <= '0;
        weight_4_12_reg <= '0;
        weight_4_13_reg <= '0;
        weight_4_14_reg <= '0;
        weight_4_15_reg <= '0;
        weight_4_16_reg <= '0;
        weight_4_17_reg <= '0;
        weight_4_18_reg <= '0;
        weight_4_19_reg <= '0;
        weight_4_20_reg <= '0;
        weight_4_21_reg <= '0;
        weight_4_22_reg <= '0;
        weight_4_23_reg <= '0;
        weight_4_24_reg <= '0;
        weight_4_25_reg <= '0;
        weight_4_26_reg <= '0;
        weight_4_27_reg <= '0;
        weight_4_28_reg <= '0;
        weight_4_29_reg <= '0;
        weight_4_30_reg <= '0;
        weight_4_31_reg <= '0;
        weight_4_32_reg <= '0;
        weight_4_33_reg <= '0;
        weight_4_34_reg <= '0;
        weight_4_35_reg <= '0;
        weight_4_36_reg <= '0;
        weight_4_37_reg <= '0;
        weight_4_38_reg <= '0;
        weight_4_39_reg <= '0;
        weight_4_40_reg <= '0;
        weight_4_41_reg <= '0;
        weight_4_42_reg <= '0;
        weight_4_43_reg <= '0;
        weight_4_44_reg <= '0;
        weight_4_45_reg <= '0;
        weight_4_46_reg <= '0;
        weight_4_47_reg <= '0;
        weight_4_48_reg <= '0;
        weight_4_49_reg <= '0;
        weight_4_50_reg <= '0;
        weight_4_51_reg <= '0;
        weight_4_52_reg <= '0;
        weight_4_53_reg <= '0;
        weight_4_54_reg <= '0;
        weight_4_55_reg <= '0;
        weight_4_56_reg <= '0;
        weight_4_57_reg <= '0;
        weight_4_58_reg <= '0;
        weight_4_59_reg <= '0;
        weight_4_60_reg <= '0;
        weight_4_61_reg <= '0;
        weight_4_62_reg <= '0;
    end else begin
        en_reg_2 <= en_reg_1;
        weight_4_0_reg <= weight_4_0;
        weight_4_1_reg <= weight_4_1;
        weight_4_2_reg <= weight_4_2;
        weight_4_3_reg <= weight_4_3;
        weight_4_4_reg <= weight_4_4;
        weight_4_5_reg <= weight_4_5;
        weight_4_6_reg <= weight_4_6;
        weight_4_7_reg <= weight_4_7;
        weight_4_8_reg <= weight_4_8;
        weight_4_9_reg <= weight_4_9;
        weight_4_10_reg <= weight_4_10;
        weight_4_11_reg <= weight_4_11;
        weight_4_12_reg <= weight_4_12;
        weight_4_13_reg <= weight_4_13;
        weight_4_14_reg <= weight_4_14;
        weight_4_15_reg <= weight_4_15;
        weight_4_16_reg <= weight_4_16;
        weight_4_17_reg <= weight_4_17;
        weight_4_18_reg <= weight_4_18;
        weight_4_19_reg <= weight_4_19;
        weight_4_20_reg <= weight_4_20;
        weight_4_21_reg <= weight_4_21;
        weight_4_22_reg <= weight_4_22;
        weight_4_23_reg <= weight_4_23;
        weight_4_24_reg <= weight_4_24;
        weight_4_25_reg <= weight_4_25;
        weight_4_26_reg <= weight_4_26;
        weight_4_27_reg <= weight_4_27;
        weight_4_28_reg <= weight_4_28;
        weight_4_29_reg <= weight_4_29;
        weight_4_30_reg <= weight_4_30;
        weight_4_31_reg <= weight_4_31;
        weight_4_32_reg <= weight_4_32;
        weight_4_33_reg <= weight_4_33;
        weight_4_34_reg <= weight_4_34;
        weight_4_35_reg <= weight_4_35;
        weight_4_36_reg <= weight_4_36;
        weight_4_37_reg <= weight_4_37;
        weight_4_38_reg <= weight_4_38;
        weight_4_39_reg <= weight_4_39;
        weight_4_40_reg <= weight_4_40;
        weight_4_41_reg <= weight_4_41;
        weight_4_42_reg <= weight_4_42;
        weight_4_43_reg <= weight_4_43;
        weight_4_44_reg <= weight_4_44;
        weight_4_45_reg <= weight_4_45;
        weight_4_46_reg <= weight_4_46;
        weight_4_47_reg <= weight_4_47;
        weight_4_48_reg <= weight_4_48;
        weight_4_49_reg <= weight_4_49;
        weight_4_50_reg <= weight_4_50;
        weight_4_51_reg <= weight_4_51;
        weight_4_52_reg <= weight_4_52;
        weight_4_53_reg <= weight_4_53;
        weight_4_54_reg <= weight_4_54;
        weight_4_55_reg <= weight_4_55;
        weight_4_56_reg <= weight_4_56;
        weight_4_57_reg <= weight_4_57;
        weight_4_58_reg <= weight_4_58;
        weight_4_59_reg <= weight_4_59;
        weight_4_60_reg <= weight_4_60;
        weight_4_61_reg <= weight_4_61;
        weight_4_62_reg <= weight_4_62;
    end
end

assign weight_4_0 = weight_3_0;
assign weight_4_1 = weight_3_1;
assign weight_4_2 = weight_3_2;
assign weight_4_3 = weight_3_3;
half_adder ha58(.a(weight_3_4[0]), .b(weight_3_4[1]), .sum(weight_4_4), .cout(weight_4_5[0]));
half_adder ha59(.a(weight_3_5[0]), .b(weight_3_5[1]), .sum(weight_4_5[1]), .cout(weight_4_6[0]));
half_adder ha60(.a(weight_3_6[0]), .b(weight_3_6[1]), .sum(weight_4_6[1]), .cout(weight_4_7[0]));
full_adder fa662(.a(weight_3_7[0]), .b(weight_3_7[1]), .cin(weight_3_7[2]), .sum(weight_4_7[1]), .cout(weight_4_8[0]));
full_adder fa663(.a(weight_3_8[0]), .b(weight_3_8[1]), .cin(weight_3_8[2]), .sum(weight_4_8[1]), .cout(weight_4_9[0]));
full_adder fa664(.a(weight_3_9[0]), .b(weight_3_9[1]), .cin(weight_3_9[2]), .sum(weight_4_9[1]), .cout(weight_4_10[0]));
full_adder fa665(.a(weight_3_10[0]), .b(weight_3_10[1]), .cin(weight_3_10[2]), .sum(weight_4_10[1]), .cout(weight_4_11[0]));
full_adder fa666(.a(weight_3_11[0]), .b(weight_3_11[1]), .cin(weight_3_11[2]), .sum(weight_4_11[1]), .cout(weight_4_12[0]));
full_adder fa667(.a(weight_3_12[0]), .b(weight_3_12[1]), .cin(weight_3_12[2]), .sum(weight_4_12[1]), .cout(weight_4_13[0]));
full_adder fa668(.a(weight_3_13[0]), .b(weight_3_13[1]), .cin(weight_3_13[2]), .sum(weight_4_13[1]), .cout(weight_4_14[0]));
full_adder fa669(.a(weight_3_14[0]), .b(weight_3_14[1]), .cin(weight_3_14[2]), .sum(weight_4_14[1]), .cout(weight_4_15[0]));
full_adder fa670(.a(weight_3_15[0]), .b(weight_3_15[1]), .cin(weight_3_15[2]), .sum(weight_4_15[1]), .cout(weight_4_16[0]));
full_adder fa671(.a(weight_3_16[0]), .b(weight_3_16[1]), .cin(weight_3_16[2]), .sum(weight_4_16[1]), .cout(weight_4_17[0]));
full_adder fa672(.a(weight_3_17[0]), .b(weight_3_17[1]), .cin(weight_3_17[2]), .sum(weight_4_17[1]), .cout(weight_4_18[0]));
full_adder fa673(.a(weight_3_18[0]), .b(weight_3_18[1]), .cin(weight_3_18[2]), .sum(weight_4_18[1]), .cout(weight_4_19[0]));
full_adder fa674(.a(weight_3_19[0]), .b(weight_3_19[1]), .cin(weight_3_19[2]), .sum(weight_4_19[1]), .cout(weight_4_20[0]));
full_adder fa675(.a(weight_3_20[0]), .b(weight_3_20[1]), .cin(weight_3_20[2]), .sum(weight_4_20[1]), .cout(weight_4_21[0]));
full_adder fa676(.a(weight_3_21[0]), .b(weight_3_21[1]), .cin(weight_3_21[2]), .sum(weight_4_21[1]), .cout(weight_4_22[0]));
full_adder fa677(.a(weight_3_22[0]), .b(weight_3_22[1]), .cin(weight_3_22[2]), .sum(weight_4_22[1]), .cout(weight_4_23[0]));
full_adder fa678(.a(weight_3_23[0]), .b(weight_3_23[1]), .cin(weight_3_23[2]), .sum(weight_4_23[1]), .cout(weight_4_24[0]));
full_adder fa679(.a(weight_3_24[0]), .b(weight_3_24[1]), .cin(weight_3_24[2]), .sum(weight_4_24[1]), .cout(weight_4_25[0]));
full_adder fa680(.a(weight_3_25[0]), .b(weight_3_25[1]), .cin(weight_3_25[2]), .sum(weight_4_25[1]), .cout(weight_4_26[0]));
full_adder fa681(.a(weight_3_26[0]), .b(weight_3_26[1]), .cin(weight_3_26[2]), .sum(weight_4_26[1]), .cout(weight_4_27[0]));
full_adder fa682(.a(weight_3_27[0]), .b(weight_3_27[1]), .cin(weight_3_27[2]), .sum(weight_4_27[1]), .cout(weight_4_28[0]));
full_adder fa683(.a(weight_3_28[0]), .b(weight_3_28[1]), .cin(weight_3_28[2]), .sum(weight_4_28[1]), .cout(weight_4_29[0]));
full_adder fa684(.a(weight_3_29[0]), .b(weight_3_29[1]), .cin(weight_3_29[2]), .sum(weight_4_29[1]), .cout(weight_4_30[0]));
full_adder fa685(.a(weight_3_30[0]), .b(weight_3_30[1]), .cin(weight_3_30[2]), .sum(weight_4_30[1]), .cout(weight_4_31[0]));
full_adder fa686(.a(weight_3_31[0]), .b(weight_3_31[1]), .cin(weight_3_31[2]), .sum(weight_4_31[1]), .cout(weight_4_32[0]));
full_adder fa687(.a(weight_3_32[0]), .b(weight_3_32[1]), .cin(weight_3_32[2]), .sum(weight_4_32[1]), .cout(weight_4_33[0]));
full_adder fa688(.a(weight_3_33[0]), .b(weight_3_33[1]), .cin(weight_3_33[2]), .sum(weight_4_33[1]), .cout(weight_4_34[0]));
full_adder fa689(.a(weight_3_34[0]), .b(weight_3_34[1]), .cin(weight_3_34[2]), .sum(weight_4_34[1]), .cout(weight_4_35[0]));
full_adder fa690(.a(weight_3_35[0]), .b(weight_3_35[1]), .cin(weight_3_35[2]), .sum(weight_4_35[1]), .cout(weight_4_36[0]));
full_adder fa691(.a(weight_3_36[0]), .b(weight_3_36[1]), .cin(weight_3_36[2]), .sum(weight_4_36[1]), .cout(weight_4_37[0]));
full_adder fa692(.a(weight_3_37[0]), .b(weight_3_37[1]), .cin(weight_3_37[2]), .sum(weight_4_37[1]), .cout(weight_4_38[0]));
half_adder ha61(.a(weight_3_38[0]), .b(weight_3_38[1]), .sum(weight_4_38[1]), .cout(weight_4_39[0]));
half_adder ha62(.a(weight_3_39[0]), .b(weight_3_39[1]), .sum(weight_4_39[1]), .cout(weight_4_40[0]));
assign weight_4_40[1] = weight_3_40[0];
assign weight_4_41[0] = weight_3_41[0];
assign weight_4_42[0] = weight_3_42[0];
assign weight_4_43[0] = weight_3_43[0];
assign weight_4_44[0] = weight_3_44[0];
assign weight_4_10[2] = weight_3_10[3];
assign weight_4_11[2] = weight_3_11[3];
assign weight_4_12[2] = weight_3_12[3];
assign weight_4_13[2] = weight_3_13[3];
half_adder ha63(.a(weight_3_14[3]), .b(weight_3_14[4]), .sum(weight_4_14[2]), .cout(weight_4_15[2]));
half_adder ha64(.a(weight_3_15[3]), .b(weight_3_15[4]), .sum(weight_4_15[3]), .cout(weight_4_16[2]));
half_adder ha65(.a(weight_3_16[3]), .b(weight_3_16[4]), .sum(weight_4_16[3]), .cout(weight_4_17[2]));
full_adder fa693(.a(weight_3_17[3]), .b(weight_3_17[4]), .cin(weight_3_17[5]), .sum(weight_4_17[3]), .cout(weight_4_18[2]));
full_adder fa694(.a(weight_3_18[3]), .b(weight_3_18[4]), .cin(weight_3_18[5]), .sum(weight_4_18[3]), .cout(weight_4_19[2]));
full_adder fa695(.a(weight_3_19[3]), .b(weight_3_19[4]), .cin(weight_3_19[5]), .sum(weight_4_19[3]), .cout(weight_4_20[2]));
full_adder fa696(.a(weight_3_20[3]), .b(weight_3_20[4]), .cin(weight_3_20[5]), .sum(weight_4_20[3]), .cout(weight_4_21[2]));
full_adder fa697(.a(weight_3_21[3]), .b(weight_3_21[4]), .cin(weight_3_21[5]), .sum(weight_4_21[3]), .cout(weight_4_22[2]));
full_adder fa698(.a(weight_3_22[3]), .b(weight_3_22[4]), .cin(weight_3_22[5]), .sum(weight_4_22[3]), .cout(weight_4_23[2]));
full_adder fa699(.a(weight_3_23[3]), .b(weight_3_23[4]), .cin(weight_3_23[5]), .sum(weight_4_23[3]), .cout(weight_4_24[2]));
full_adder fa700(.a(weight_3_24[3]), .b(weight_3_24[4]), .cin(weight_3_24[5]), .sum(weight_4_24[3]), .cout(weight_4_25[2]));
full_adder fa701(.a(weight_3_25[3]), .b(weight_3_25[4]), .cin(weight_3_25[5]), .sum(weight_4_25[3]), .cout(weight_4_26[2]));
full_adder fa702(.a(weight_3_26[3]), .b(weight_3_26[4]), .cin(weight_3_26[5]), .sum(weight_4_26[3]), .cout(weight_4_27[2]));
full_adder fa703(.a(weight_3_27[3]), .b(weight_3_27[4]), .cin(weight_3_27[5]), .sum(weight_4_27[3]), .cout(weight_4_28[2]));
full_adder fa704(.a(weight_3_28[3]), .b(weight_3_28[4]), .cin(weight_3_28[5]), .sum(weight_4_28[3]), .cout(weight_4_29[2]));
full_adder fa705(.a(weight_3_29[3]), .b(weight_3_29[4]), .cin(weight_3_29[5]), .sum(weight_4_29[3]), .cout(weight_4_30[2]));
full_adder fa706(.a(weight_3_30[3]), .b(weight_3_30[4]), .cin(weight_3_30[5]), .sum(weight_4_30[3]), .cout(weight_4_31[2]));
full_adder fa707(.a(weight_3_31[3]), .b(weight_3_31[4]), .cin(weight_3_31[5]), .sum(weight_4_31[3]), .cout(weight_4_32[2]));
full_adder fa708(.a(weight_3_32[3]), .b(weight_3_32[4]), .cin(weight_3_32[5]), .sum(weight_4_32[3]), .cout(weight_4_33[2]));
full_adder fa709(.a(weight_3_33[3]), .b(weight_3_33[4]), .cin(weight_3_33[5]), .sum(weight_4_33[3]), .cout(weight_4_34[2]));
full_adder fa710(.a(weight_3_34[3]), .b(weight_3_34[4]), .cin(weight_3_34[5]), .sum(weight_4_34[3]), .cout(weight_4_35[2]));
full_adder fa711(.a(weight_3_35[3]), .b(weight_3_35[4]), .cin(weight_3_35[5]), .sum(weight_4_35[3]), .cout(weight_4_36[2]));
full_adder fa712(.a(weight_3_36[3]), .b(weight_3_36[4]), .cin(weight_3_36[5]), .sum(weight_4_36[3]), .cout(weight_4_37[2]));
full_adder fa713(.a(weight_3_37[3]), .b(weight_3_37[4]), .cin(weight_3_37[5]), .sum(weight_4_37[3]), .cout(weight_4_38[2]));
full_adder fa714(.a(weight_3_38[2]), .b(weight_3_38[3]), .cin(weight_3_38[4]), .sum(weight_4_38[3]), .cout(weight_4_39[2]));
full_adder fa715(.a(weight_3_39[2]), .b(weight_3_39[3]), .cin(weight_3_39[4]), .sum(weight_4_39[3]), .cout(weight_4_40[2]));
full_adder fa716(.a(weight_3_40[1]), .b(weight_3_40[2]), .cin(weight_3_40[3]), .sum(weight_4_40[3]), .cout(weight_4_41[1]));
full_adder fa717(.a(weight_3_41[1]), .b(weight_3_41[2]), .cin(weight_3_41[3]), .sum(weight_4_41[2]), .cout(weight_4_42[1]));
full_adder fa718(.a(weight_3_42[1]), .b(weight_3_42[2]), .cin(weight_3_42[3]), .sum(weight_4_42[2]), .cout(weight_4_43[1]));
full_adder fa719(.a(weight_3_43[1]), .b(weight_3_43[2]), .cin(weight_3_43[3]), .sum(weight_4_43[2]), .cout(weight_4_44[1]));
full_adder fa720(.a(weight_3_44[1]), .b(weight_3_44[2]), .cin(weight_3_44[3]), .sum(weight_4_44[2]), .cout(weight_4_45[0]));
full_adder fa721(.a(weight_3_45[0]), .b(weight_3_45[1]), .cin(weight_3_45[2]), .sum(weight_4_45[1]), .cout(weight_4_46[0]));
half_adder ha66(.a(weight_3_46[0]), .b(weight_3_46[1]), .sum(weight_4_46[1]), .cout(weight_4_47[0]));
half_adder ha67(.a(weight_3_47[0]), .b(weight_3_47[1]), .sum(weight_4_47[1]), .cout(weight_4_48[0]));
half_adder ha68(.a(weight_3_48[0]), .b(weight_3_48[1]), .sum(weight_4_48[1]), .cout(weight_4_49[0]));
half_adder ha69(.a(weight_3_49[0]), .b(weight_3_49[1]), .sum(weight_4_49[1]), .cout(weight_4_50[0]));
half_adder ha70(.a(weight_3_50[0]), .b(weight_3_50[1]), .sum(weight_4_50[1]), .cout(weight_4_51[0]));
assign weight_4_51[1] = weight_3_51[0];
assign weight_4_52[0] = weight_3_52[0];
assign weight_4_21[4] = weight_3_21[6];
assign weight_4_22[4] = weight_3_22[6];
assign weight_4_23[4] = weight_3_23[6];
half_adder ha71(.a(weight_3_24[6]), .b(weight_3_24[7]), .sum(weight_4_24[4]), .cout(weight_4_25[4]));
half_adder ha72(.a(weight_3_25[6]), .b(weight_3_25[7]), .sum(weight_4_25[5]), .cout(weight_4_26[4]));
half_adder ha73(.a(weight_3_26[6]), .b(weight_3_26[7]), .sum(weight_4_26[5]), .cout(weight_4_27[4]));
full_adder fa722(.a(weight_3_27[6]), .b(weight_3_27[7]), .cin(weight_3_27[8]), .sum(weight_4_27[5]), .cout(weight_4_28[4]));
full_adder fa723(.a(weight_3_28[6]), .b(weight_3_28[7]), .cin(weight_3_28[8]), .sum(weight_4_28[5]), .cout(weight_4_29[4]));
full_adder fa724(.a(weight_3_29[6]), .b(weight_3_29[7]), .cin(weight_3_29[8]), .sum(weight_4_29[5]), .cout(weight_4_30[4]));
full_adder fa725(.a(weight_3_30[6]), .b(weight_3_30[7]), .cin(weight_3_30[8]), .sum(weight_4_30[5]), .cout(weight_4_31[4]));
full_adder fa726(.a(weight_3_31[6]), .b(weight_3_31[7]), .cin(weight_3_31[8]), .sum(weight_4_31[5]), .cout(weight_4_32[4]));
full_adder fa727(.a(weight_3_32[6]), .b(weight_3_32[7]), .cin(weight_3_32[8]), .sum(weight_4_32[5]), .cout(weight_4_33[4]));
full_adder fa728(.a(weight_3_33[6]), .b(weight_3_33[7]), .cin(weight_3_33[8]), .sum(weight_4_33[5]), .cout(weight_4_34[4]));
full_adder fa729(.a(weight_3_34[6]), .b(weight_3_34[7]), .cin(weight_3_34[8]), .sum(weight_4_34[5]), .cout(weight_4_35[4]));
full_adder fa730(.a(weight_3_35[6]), .b(weight_3_35[7]), .cin(weight_3_35[8]), .sum(weight_4_35[5]), .cout(weight_4_36[4]));
full_adder fa731(.a(weight_3_36[6]), .b(weight_3_36[7]), .cin(weight_3_36[8]), .sum(weight_4_36[5]), .cout(weight_4_37[4]));
full_adder fa732(.a(weight_3_37[6]), .b(weight_3_37[7]), .cin(weight_3_37[8]), .sum(weight_4_37[5]), .cout(weight_4_38[4]));
full_adder fa733(.a(weight_3_38[5]), .b(weight_3_38[6]), .cin(weight_3_38[7]), .sum(weight_4_38[5]), .cout(weight_4_39[4]));
full_adder fa734(.a(weight_3_39[5]), .b(weight_3_39[6]), .cin(weight_3_39[7]), .sum(weight_4_39[5]), .cout(weight_4_40[4]));
full_adder fa735(.a(weight_3_40[4]), .b(weight_3_40[5]), .cin(weight_3_40[6]), .sum(weight_4_40[5]), .cout(weight_4_41[3]));
full_adder fa736(.a(weight_3_41[4]), .b(weight_3_41[5]), .cin(weight_3_41[6]), .sum(weight_4_41[4]), .cout(weight_4_42[3]));
full_adder fa737(.a(weight_3_42[4]), .b(weight_3_42[5]), .cin(weight_3_42[6]), .sum(weight_4_42[4]), .cout(weight_4_43[3]));
full_adder fa738(.a(weight_3_43[4]), .b(weight_3_43[5]), .cin(weight_3_43[6]), .sum(weight_4_43[4]), .cout(weight_4_44[3]));
full_adder fa739(.a(weight_3_44[4]), .b(weight_3_44[5]), .cin(weight_3_44[6]), .sum(weight_4_44[4]), .cout(weight_4_45[2]));
full_adder fa740(.a(weight_3_45[3]), .b(weight_3_45[4]), .cin(weight_3_45[5]), .sum(weight_4_45[3]), .cout(weight_4_46[2]));
full_adder fa741(.a(weight_3_46[2]), .b(weight_3_46[3]), .cin(weight_3_46[4]), .sum(weight_4_46[3]), .cout(weight_4_47[2]));
full_adder fa742(.a(weight_3_47[2]), .b(weight_3_47[3]), .cin(weight_3_47[4]), .sum(weight_4_47[3]), .cout(weight_4_48[2]));
full_adder fa743(.a(weight_3_48[2]), .b(weight_3_48[3]), .cin(weight_3_48[4]), .sum(weight_4_48[3]), .cout(weight_4_49[2]));
full_adder fa744(.a(weight_3_49[2]), .b(weight_3_49[3]), .cin(weight_3_49[4]), .sum(weight_4_49[3]), .cout(weight_4_50[2]));
full_adder fa745(.a(weight_3_50[2]), .b(weight_3_50[3]), .cin(weight_3_50[4]), .sum(weight_4_50[3]), .cout(weight_4_51[2]));
full_adder fa746(.a(weight_3_51[1]), .b(weight_3_51[2]), .cin(weight_3_51[3]), .sum(weight_4_51[3]), .cout(weight_4_52[1]));
full_adder fa747(.a(weight_3_52[1]), .b(weight_3_52[2]), .cin(weight_3_52[3]), .sum(weight_4_52[2]), .cout(weight_4_53[0]));
full_adder fa748(.a(weight_3_53[0]), .b(weight_3_53[1]), .cin(weight_3_53[2]), .sum(weight_4_53[1]), .cout(weight_4_54[0]));
full_adder fa749(.a(weight_3_54[0]), .b(weight_3_54[1]), .cin(weight_3_54[2]), .sum(weight_4_54[1]), .cout(weight_4_55[0]));
full_adder fa750(.a(weight_3_55[0]), .b(weight_3_55[1]), .cin(weight_3_55[2]), .sum(weight_4_55[1]), .cout(weight_4_56[0]));
full_adder fa751(.a(weight_3_56[0]), .b(weight_3_56[1]), .cin(weight_3_56[2]), .sum(weight_4_56[1]), .cout(weight_4_57[0]));
full_adder fa752(.a(weight_3_57[0]), .b(weight_3_57[1]), .cin(weight_3_57[2]), .sum(weight_4_57[1]), .cout(weight_4_58[0]));
full_adder fa753(.a(weight_3_58[0]), .b(weight_3_58[1]), .cin(weight_3_58[2]), .sum(weight_4_58[1]), .cout(weight_4_59[0]));
assign weight_4_59[1] = weight_3_59[0];
assign weight_4_60[0] = weight_3_60[0];
assign weight_4_61[0] = weight_3_61[0];
assign weight_4_62[0] = weight_3_62[0];
assign weight_4_31[6] = weight_3_31[9];
assign weight_4_32[6] = weight_3_32[9];
assign weight_4_33[6] = weight_3_33[9];
assign weight_4_34[6] = weight_3_34[9];
assign weight_4_35[6] = weight_3_35[9];
assign weight_4_36[6] = weight_3_36[9];
assign weight_4_37[6] = weight_3_37[9];
assign weight_4_38[6] = weight_3_38[8];
assign weight_4_39[6] = weight_3_39[8];
assign weight_4_40[6] = weight_3_40[7];
assign weight_4_41[5] = weight_3_41[7];
assign weight_4_42[5] = weight_3_42[7];
assign weight_4_43[5] = weight_3_43[7];
assign weight_4_44[5] = weight_3_44[7];
assign weight_4_45[4] = weight_3_45[6];
assign weight_4_46[4] = weight_3_46[5];
assign weight_4_47[4] = weight_3_47[5];
assign weight_4_48[4] = weight_3_48[5];
assign weight_4_49[4] = weight_3_49[5];
assign weight_4_50[4] = weight_3_50[5];
assign weight_4_51[4] = weight_3_51[4];
assign weight_4_52[3] = weight_3_52[4];
assign weight_4_53[2] = weight_3_53[3];
assign weight_4_54[2] = weight_3_54[3];
assign weight_4_55[2] = weight_3_55[3];
assign weight_4_56[2] = weight_3_56[3];
assign weight_4_57[2] = weight_3_57[3];
assign weight_4_58[2] = weight_3_58[3];
assign weight_4_59[2] = weight_3_59[1];
assign weight_4_60[1] = weight_3_60[1];
assign weight_4_61[1] = weight_3_61[1];
assign weight_4_62[1] = weight_3_62[1];
logic weight_5_0;
logic weight_5_1;
logic weight_5_2;
logic weight_5_3;
logic weight_5_4;
logic weight_5_5;
logic [1:0] weight_5_6;
logic [1:0] weight_5_7;
logic [1:0] weight_5_8;
logic [1:0] weight_5_9;
logic [1:0] weight_5_10;
logic [1:0] weight_5_11;
logic [1:0] weight_5_12;
logic [1:0] weight_5_13;
logic [1:0] weight_5_14;
logic [2:0] weight_5_15;
logic [2:0] weight_5_16;
logic [2:0] weight_5_17;
logic [2:0] weight_5_18;
logic [2:0] weight_5_19;
logic [2:0] weight_5_20;
logic [2:0] weight_5_21;
logic [3:0] weight_5_22;
logic [3:0] weight_5_23;
logic [3:0] weight_5_24;
logic [3:0] weight_5_25;
logic [3:0] weight_5_26;
logic [3:0] weight_5_27;
logic [3:0] weight_5_28;
logic [3:0] weight_5_29;
logic [3:0] weight_5_30;
logic [4:0] weight_5_31;
logic [4:0] weight_5_32;
logic [4:0] weight_5_33;
logic [4:0] weight_5_34;
logic [4:0] weight_5_35;
logic [4:0] weight_5_36;
logic [4:0] weight_5_37;
logic [4:0] weight_5_38;
logic [4:0] weight_5_39;
logic [4:0] weight_5_40;
logic [4:0] weight_5_41;
logic [4:0] weight_5_42;
logic [4:0] weight_5_43;
logic [4:0] weight_5_44;
logic [4:0] weight_5_45;
logic [3:0] weight_5_46;
logic [3:0] weight_5_47;
logic [3:0] weight_5_48;
logic [3:0] weight_5_49;
logic [3:0] weight_5_50;
logic [3:0] weight_5_51;
logic [2:0] weight_5_52;
logic [2:0] weight_5_53;
logic [2:0] weight_5_54;
logic [2:0] weight_5_55;
logic [2:0] weight_5_56;
logic [2:0] weight_5_57;
logic [2:0] weight_5_58;
logic [2:0] weight_5_59;
logic [2:0] weight_5_60;
logic [1:0] weight_5_61;
logic [1:0] weight_5_62;
assign weight_5_0 = weight_4_0_reg;
assign weight_5_1 = weight_4_1_reg;
assign weight_5_2 = weight_4_2_reg;
assign weight_5_3 = weight_4_3_reg;
assign weight_5_4 = weight_4_4_reg;
half_adder ha74(.a(weight_4_5_reg[0]), .b(weight_4_5_reg[1]), .sum(weight_5_5), .cout(weight_5_6[0]));
half_adder ha75(.a(weight_4_6_reg[0]), .b(weight_4_6_reg[1]), .sum(weight_5_6[1]), .cout(weight_5_7[0]));
half_adder ha76(.a(weight_4_7_reg[0]), .b(weight_4_7_reg[1]), .sum(weight_5_7[1]), .cout(weight_5_8[0]));
half_adder ha77(.a(weight_4_8_reg[0]), .b(weight_4_8_reg[1]), .sum(weight_5_8[1]), .cout(weight_5_9[0]));
half_adder ha78(.a(weight_4_9_reg[0]), .b(weight_4_9_reg[1]), .sum(weight_5_9[1]), .cout(weight_5_10[0]));
full_adder fa754(.a(weight_4_10_reg[0]), .b(weight_4_10_reg[1]), .cin(weight_4_10_reg[2]), .sum(weight_5_10[1]), .cout(weight_5_11[0]));
full_adder fa755(.a(weight_4_11_reg[0]), .b(weight_4_11_reg[1]), .cin(weight_4_11_reg[2]), .sum(weight_5_11[1]), .cout(weight_5_12[0]));
full_adder fa756(.a(weight_4_12_reg[0]), .b(weight_4_12_reg[1]), .cin(weight_4_12_reg[2]), .sum(weight_5_12[1]), .cout(weight_5_13[0]));
full_adder fa757(.a(weight_4_13_reg[0]), .b(weight_4_13_reg[1]), .cin(weight_4_13_reg[2]), .sum(weight_5_13[1]), .cout(weight_5_14[0]));
full_adder fa758(.a(weight_4_14_reg[0]), .b(weight_4_14_reg[1]), .cin(weight_4_14_reg[2]), .sum(weight_5_14[1]), .cout(weight_5_15[0]));
full_adder fa759(.a(weight_4_15_reg[0]), .b(weight_4_15_reg[1]), .cin(weight_4_15_reg[2]), .sum(weight_5_15[1]), .cout(weight_5_16[0]));
full_adder fa760(.a(weight_4_16_reg[0]), .b(weight_4_16_reg[1]), .cin(weight_4_16_reg[2]), .sum(weight_5_16[1]), .cout(weight_5_17[0]));
full_adder fa761(.a(weight_4_17_reg[0]), .b(weight_4_17_reg[1]), .cin(weight_4_17_reg[2]), .sum(weight_5_17[1]), .cout(weight_5_18[0]));
full_adder fa762(.a(weight_4_18_reg[0]), .b(weight_4_18_reg[1]), .cin(weight_4_18_reg[2]), .sum(weight_5_18[1]), .cout(weight_5_19[0]));
full_adder fa763(.a(weight_4_19_reg[0]), .b(weight_4_19_reg[1]), .cin(weight_4_19_reg[2]), .sum(weight_5_19[1]), .cout(weight_5_20[0]));
full_adder fa764(.a(weight_4_20_reg[0]), .b(weight_4_20_reg[1]), .cin(weight_4_20_reg[2]), .sum(weight_5_20[1]), .cout(weight_5_21[0]));
full_adder fa765(.a(weight_4_21_reg[0]), .b(weight_4_21_reg[1]), .cin(weight_4_21_reg[2]), .sum(weight_5_21[1]), .cout(weight_5_22[0]));
full_adder fa766(.a(weight_4_22_reg[0]), .b(weight_4_22_reg[1]), .cin(weight_4_22_reg[2]), .sum(weight_5_22[1]), .cout(weight_5_23[0]));
full_adder fa767(.a(weight_4_23_reg[0]), .b(weight_4_23_reg[1]), .cin(weight_4_23_reg[2]), .sum(weight_5_23[1]), .cout(weight_5_24[0]));
full_adder fa768(.a(weight_4_24_reg[0]), .b(weight_4_24_reg[1]), .cin(weight_4_24_reg[2]), .sum(weight_5_24[1]), .cout(weight_5_25[0]));
full_adder fa769(.a(weight_4_25_reg[0]), .b(weight_4_25_reg[1]), .cin(weight_4_25_reg[2]), .sum(weight_5_25[1]), .cout(weight_5_26[0]));
full_adder fa770(.a(weight_4_26_reg[0]), .b(weight_4_26_reg[1]), .cin(weight_4_26_reg[2]), .sum(weight_5_26[1]), .cout(weight_5_27[0]));
full_adder fa771(.a(weight_4_27_reg[0]), .b(weight_4_27_reg[1]), .cin(weight_4_27_reg[2]), .sum(weight_5_27[1]), .cout(weight_5_28[0]));
full_adder fa772(.a(weight_4_28_reg[0]), .b(weight_4_28_reg[1]), .cin(weight_4_28_reg[2]), .sum(weight_5_28[1]), .cout(weight_5_29[0]));
full_adder fa773(.a(weight_4_29_reg[0]), .b(weight_4_29_reg[1]), .cin(weight_4_29_reg[2]), .sum(weight_5_29[1]), .cout(weight_5_30[0]));
full_adder fa774(.a(weight_4_30_reg[0]), .b(weight_4_30_reg[1]), .cin(weight_4_30_reg[2]), .sum(weight_5_30[1]), .cout(weight_5_31[0]));
full_adder fa775(.a(weight_4_31_reg[0]), .b(weight_4_31_reg[1]), .cin(weight_4_31_reg[2]), .sum(weight_5_31[1]), .cout(weight_5_32[0]));
full_adder fa776(.a(weight_4_32_reg[0]), .b(weight_4_32_reg[1]), .cin(weight_4_32_reg[2]), .sum(weight_5_32[1]), .cout(weight_5_33[0]));
full_adder fa777(.a(weight_4_33_reg[0]), .b(weight_4_33_reg[1]), .cin(weight_4_33_reg[2]), .sum(weight_5_33[1]), .cout(weight_5_34[0]));
full_adder fa778(.a(weight_4_34_reg[0]), .b(weight_4_34_reg[1]), .cin(weight_4_34_reg[2]), .sum(weight_5_34[1]), .cout(weight_5_35[0]));
full_adder fa779(.a(weight_4_35_reg[0]), .b(weight_4_35_reg[1]), .cin(weight_4_35_reg[2]), .sum(weight_5_35[1]), .cout(weight_5_36[0]));
full_adder fa780(.a(weight_4_36_reg[0]), .b(weight_4_36_reg[1]), .cin(weight_4_36_reg[2]), .sum(weight_5_36[1]), .cout(weight_5_37[0]));
full_adder fa781(.a(weight_4_37_reg[0]), .b(weight_4_37_reg[1]), .cin(weight_4_37_reg[2]), .sum(weight_5_37[1]), .cout(weight_5_38[0]));
full_adder fa782(.a(weight_4_38_reg[0]), .b(weight_4_38_reg[1]), .cin(weight_4_38_reg[2]), .sum(weight_5_38[1]), .cout(weight_5_39[0]));
full_adder fa783(.a(weight_4_39_reg[0]), .b(weight_4_39_reg[1]), .cin(weight_4_39_reg[2]), .sum(weight_5_39[1]), .cout(weight_5_40[0]));
full_adder fa784(.a(weight_4_40_reg[0]), .b(weight_4_40_reg[1]), .cin(weight_4_40_reg[2]), .sum(weight_5_40[1]), .cout(weight_5_41[0]));
half_adder ha79(.a(weight_4_41_reg[0]), .b(weight_4_41_reg[1]), .sum(weight_5_41[1]), .cout(weight_5_42[0]));
half_adder ha80(.a(weight_4_42_reg[0]), .b(weight_4_42_reg[1]), .sum(weight_5_42[1]), .cout(weight_5_43[0]));
half_adder ha81(.a(weight_4_43_reg[0]), .b(weight_4_43_reg[1]), .sum(weight_5_43[1]), .cout(weight_5_44[0]));
half_adder ha82(.a(weight_4_44_reg[0]), .b(weight_4_44_reg[1]), .sum(weight_5_44[1]), .cout(weight_5_45[0]));
assign weight_5_45[1] = weight_4_45_reg[0];
assign weight_5_46[0] = weight_4_46_reg[0];
assign weight_5_47[0] = weight_4_47_reg[0];
assign weight_5_48[0] = weight_4_48_reg[0];
assign weight_5_49[0] = weight_4_49_reg[0];
assign weight_5_50[0] = weight_4_50_reg[0];
assign weight_5_51[0] = weight_4_51_reg[0];
assign weight_5_15[2] = weight_4_15_reg[3];
assign weight_5_16[2] = weight_4_16_reg[3];
assign weight_5_17[2] = weight_4_17_reg[3];
assign weight_5_18[2] = weight_4_18_reg[3];
assign weight_5_19[2] = weight_4_19_reg[3];
assign weight_5_20[2] = weight_4_20_reg[3];
half_adder ha83(.a(weight_4_21_reg[3]), .b(weight_4_21_reg[4]), .sum(weight_5_21[2]), .cout(weight_5_22[2]));
half_adder ha84(.a(weight_4_22_reg[3]), .b(weight_4_22_reg[4]), .sum(weight_5_22[3]), .cout(weight_5_23[2]));
half_adder ha85(.a(weight_4_23_reg[3]), .b(weight_4_23_reg[4]), .sum(weight_5_23[3]), .cout(weight_5_24[2]));
half_adder ha86(.a(weight_4_24_reg[3]), .b(weight_4_24_reg[4]), .sum(weight_5_24[3]), .cout(weight_5_25[2]));
full_adder fa785(.a(weight_4_25_reg[3]), .b(weight_4_25_reg[4]), .cin(weight_4_25_reg[5]), .sum(weight_5_25[3]), .cout(weight_5_26[2]));
full_adder fa786(.a(weight_4_26_reg[3]), .b(weight_4_26_reg[4]), .cin(weight_4_26_reg[5]), .sum(weight_5_26[3]), .cout(weight_5_27[2]));
full_adder fa787(.a(weight_4_27_reg[3]), .b(weight_4_27_reg[4]), .cin(weight_4_27_reg[5]), .sum(weight_5_27[3]), .cout(weight_5_28[2]));
full_adder fa788(.a(weight_4_28_reg[3]), .b(weight_4_28_reg[4]), .cin(weight_4_28_reg[5]), .sum(weight_5_28[3]), .cout(weight_5_29[2]));
full_adder fa789(.a(weight_4_29_reg[3]), .b(weight_4_29_reg[4]), .cin(weight_4_29_reg[5]), .sum(weight_5_29[3]), .cout(weight_5_30[2]));
full_adder fa790(.a(weight_4_30_reg[3]), .b(weight_4_30_reg[4]), .cin(weight_4_30_reg[5]), .sum(weight_5_30[3]), .cout(weight_5_31[2]));
full_adder fa791(.a(weight_4_31_reg[3]), .b(weight_4_31_reg[4]), .cin(weight_4_31_reg[5]), .sum(weight_5_31[3]), .cout(weight_5_32[2]));
full_adder fa792(.a(weight_4_32_reg[3]), .b(weight_4_32_reg[4]), .cin(weight_4_32_reg[5]), .sum(weight_5_32[3]), .cout(weight_5_33[2]));
full_adder fa793(.a(weight_4_33_reg[3]), .b(weight_4_33_reg[4]), .cin(weight_4_33_reg[5]), .sum(weight_5_33[3]), .cout(weight_5_34[2]));
full_adder fa794(.a(weight_4_34_reg[3]), .b(weight_4_34_reg[4]), .cin(weight_4_34_reg[5]), .sum(weight_5_34[3]), .cout(weight_5_35[2]));
full_adder fa795(.a(weight_4_35_reg[3]), .b(weight_4_35_reg[4]), .cin(weight_4_35_reg[5]), .sum(weight_5_35[3]), .cout(weight_5_36[2]));
full_adder fa796(.a(weight_4_36_reg[3]), .b(weight_4_36_reg[4]), .cin(weight_4_36_reg[5]), .sum(weight_5_36[3]), .cout(weight_5_37[2]));
full_adder fa797(.a(weight_4_37_reg[3]), .b(weight_4_37_reg[4]), .cin(weight_4_37_reg[5]), .sum(weight_5_37[3]), .cout(weight_5_38[2]));
full_adder fa798(.a(weight_4_38_reg[3]), .b(weight_4_38_reg[4]), .cin(weight_4_38_reg[5]), .sum(weight_5_38[3]), .cout(weight_5_39[2]));
full_adder fa799(.a(weight_4_39_reg[3]), .b(weight_4_39_reg[4]), .cin(weight_4_39_reg[5]), .sum(weight_5_39[3]), .cout(weight_5_40[2]));
full_adder fa800(.a(weight_4_40_reg[3]), .b(weight_4_40_reg[4]), .cin(weight_4_40_reg[5]), .sum(weight_5_40[3]), .cout(weight_5_41[2]));
full_adder fa801(.a(weight_4_41_reg[2]), .b(weight_4_41_reg[3]), .cin(weight_4_41_reg[4]), .sum(weight_5_41[3]), .cout(weight_5_42[2]));
full_adder fa802(.a(weight_4_42_reg[2]), .b(weight_4_42_reg[3]), .cin(weight_4_42_reg[4]), .sum(weight_5_42[3]), .cout(weight_5_43[2]));
full_adder fa803(.a(weight_4_43_reg[2]), .b(weight_4_43_reg[3]), .cin(weight_4_43_reg[4]), .sum(weight_5_43[3]), .cout(weight_5_44[2]));
full_adder fa804(.a(weight_4_44_reg[2]), .b(weight_4_44_reg[3]), .cin(weight_4_44_reg[4]), .sum(weight_5_44[3]), .cout(weight_5_45[2]));
full_adder fa805(.a(weight_4_45_reg[1]), .b(weight_4_45_reg[2]), .cin(weight_4_45_reg[3]), .sum(weight_5_45[3]), .cout(weight_5_46[1]));
full_adder fa806(.a(weight_4_46_reg[1]), .b(weight_4_46_reg[2]), .cin(weight_4_46_reg[3]), .sum(weight_5_46[2]), .cout(weight_5_47[1]));
full_adder fa807(.a(weight_4_47_reg[1]), .b(weight_4_47_reg[2]), .cin(weight_4_47_reg[3]), .sum(weight_5_47[2]), .cout(weight_5_48[1]));
full_adder fa808(.a(weight_4_48_reg[1]), .b(weight_4_48_reg[2]), .cin(weight_4_48_reg[3]), .sum(weight_5_48[2]), .cout(weight_5_49[1]));
full_adder fa809(.a(weight_4_49_reg[1]), .b(weight_4_49_reg[2]), .cin(weight_4_49_reg[3]), .sum(weight_5_49[2]), .cout(weight_5_50[1]));
full_adder fa810(.a(weight_4_50_reg[1]), .b(weight_4_50_reg[2]), .cin(weight_4_50_reg[3]), .sum(weight_5_50[2]), .cout(weight_5_51[1]));
full_adder fa811(.a(weight_4_51_reg[1]), .b(weight_4_51_reg[2]), .cin(weight_4_51_reg[3]), .sum(weight_5_51[2]), .cout(weight_5_52[0]));
full_adder fa812(.a(weight_4_52_reg[0]), .b(weight_4_52_reg[1]), .cin(weight_4_52_reg[2]), .sum(weight_5_52[1]), .cout(weight_5_53[0]));
half_adder ha87(.a(weight_4_53_reg[0]), .b(weight_4_53_reg[1]), .sum(weight_5_53[1]), .cout(weight_5_54[0]));
half_adder ha88(.a(weight_4_54_reg[0]), .b(weight_4_54_reg[1]), .sum(weight_5_54[1]), .cout(weight_5_55[0]));
half_adder ha89(.a(weight_4_55_reg[0]), .b(weight_4_55_reg[1]), .sum(weight_5_55[1]), .cout(weight_5_56[0]));
half_adder ha90(.a(weight_4_56_reg[0]), .b(weight_4_56_reg[1]), .sum(weight_5_56[1]), .cout(weight_5_57[0]));
half_adder ha91(.a(weight_4_57_reg[0]), .b(weight_4_57_reg[1]), .sum(weight_5_57[1]), .cout(weight_5_58[0]));
half_adder ha92(.a(weight_4_58_reg[0]), .b(weight_4_58_reg[1]), .sum(weight_5_58[1]), .cout(weight_5_59[0]));
half_adder ha93(.a(weight_4_59_reg[0]), .b(weight_4_59_reg[1]), .sum(weight_5_59[1]), .cout(weight_5_60[0]));
assign weight_5_60[1] = weight_4_60_reg[0];
assign weight_5_61[0] = weight_4_61_reg[0];
assign weight_5_62[0] = weight_4_62_reg[0];
assign weight_5_31[4] = weight_4_31_reg[6];
assign weight_5_32[4] = weight_4_32_reg[6];
assign weight_5_33[4] = weight_4_33_reg[6];
assign weight_5_34[4] = weight_4_34_reg[6];
assign weight_5_35[4] = weight_4_35_reg[6];
assign weight_5_36[4] = weight_4_36_reg[6];
assign weight_5_37[4] = weight_4_37_reg[6];
assign weight_5_38[4] = weight_4_38_reg[6];
assign weight_5_39[4] = weight_4_39_reg[6];
assign weight_5_40[4] = weight_4_40_reg[6];
assign weight_5_41[4] = weight_4_41_reg[5];
assign weight_5_42[4] = weight_4_42_reg[5];
assign weight_5_43[4] = weight_4_43_reg[5];
assign weight_5_44[4] = weight_4_44_reg[5];
assign weight_5_45[4] = weight_4_45_reg[4];
assign weight_5_46[3] = weight_4_46_reg[4];
assign weight_5_47[3] = weight_4_47_reg[4];
assign weight_5_48[3] = weight_4_48_reg[4];
assign weight_5_49[3] = weight_4_49_reg[4];
assign weight_5_50[3] = weight_4_50_reg[4];
assign weight_5_51[3] = weight_4_51_reg[4];
assign weight_5_52[2] = weight_4_52_reg[3];
assign weight_5_53[2] = weight_4_53_reg[2];
assign weight_5_54[2] = weight_4_54_reg[2];
assign weight_5_55[2] = weight_4_55_reg[2];
assign weight_5_56[2] = weight_4_56_reg[2];
assign weight_5_57[2] = weight_4_57_reg[2];
assign weight_5_58[2] = weight_4_58_reg[2];
assign weight_5_59[2] = weight_4_59_reg[2];
assign weight_5_60[2] = weight_4_60_reg[1];
assign weight_5_61[1] = weight_4_61_reg[1];
assign weight_5_62[1] = weight_4_62_reg[1];
logic weight_6_0;
logic weight_6_1;
logic weight_6_2;
logic weight_6_3;
logic weight_6_4;
logic weight_6_5;
logic weight_6_6;
logic [1:0] weight_6_7;
logic [1:0] weight_6_8;
logic [1:0] weight_6_9;
logic [1:0] weight_6_10;
logic [1:0] weight_6_11;
logic [1:0] weight_6_12;
logic [1:0] weight_6_13;
logic [1:0] weight_6_14;
logic [1:0] weight_6_15;
logic [1:0] weight_6_16;
logic [1:0] weight_6_17;
logic [1:0] weight_6_18;
logic [1:0] weight_6_19;
logic [1:0] weight_6_20;
logic [1:0] weight_6_21;
logic [2:0] weight_6_22;
logic [2:0] weight_6_23;
logic [2:0] weight_6_24;
logic [2:0] weight_6_25;
logic [2:0] weight_6_26;
logic [2:0] weight_6_27;
logic [2:0] weight_6_28;
logic [2:0] weight_6_29;
logic [2:0] weight_6_30;
logic [3:0] weight_6_31;
logic [3:0] weight_6_32;
logic [3:0] weight_6_33;
logic [3:0] weight_6_34;
logic [3:0] weight_6_35;
logic [3:0] weight_6_36;
logic [3:0] weight_6_37;
logic [3:0] weight_6_38;
logic [3:0] weight_6_39;
logic [3:0] weight_6_40;
logic [3:0] weight_6_41;
logic [3:0] weight_6_42;
logic [3:0] weight_6_43;
logic [3:0] weight_6_44;
logic [3:0] weight_6_45;
logic [3:0] weight_6_46;
logic [3:0] weight_6_47;
logic [3:0] weight_6_48;
logic [3:0] weight_6_49;
logic [3:0] weight_6_50;
logic [3:0] weight_6_51;
logic [3:0] weight_6_52;
logic [2:0] weight_6_53;
logic [2:0] weight_6_54;
logic [2:0] weight_6_55;
logic [2:0] weight_6_56;
logic [2:0] weight_6_57;
logic [2:0] weight_6_58;
logic [2:0] weight_6_59;
logic [2:0] weight_6_60;
logic [1:0] weight_6_61;
logic [1:0] weight_6_62;

logic en_reg_3;
logic weight_6_0_reg;
logic weight_6_1_reg;
logic weight_6_2_reg;
logic weight_6_3_reg;
logic weight_6_4_reg;
logic weight_6_5_reg;
logic weight_6_6_reg;
logic [1:0] weight_6_7_reg;
logic [1:0] weight_6_8_reg;
logic [1:0] weight_6_9_reg;
logic [1:0] weight_6_10_reg;
logic [1:0] weight_6_11_reg;
logic [1:0] weight_6_12_reg;
logic [1:0] weight_6_13_reg;
logic [1:0] weight_6_14_reg;
logic [1:0] weight_6_15_reg;
logic [1:0] weight_6_16_reg;
logic [1:0] weight_6_17_reg;
logic [1:0] weight_6_18_reg;
logic [1:0] weight_6_19_reg;
logic [1:0] weight_6_20_reg;
logic [1:0] weight_6_21_reg;
logic [2:0] weight_6_22_reg;
logic [2:0] weight_6_23_reg;
logic [2:0] weight_6_24_reg;
logic [2:0] weight_6_25_reg;
logic [2:0] weight_6_26_reg;
logic [2:0] weight_6_27_reg;
logic [2:0] weight_6_28_reg;
logic [2:0] weight_6_29_reg;
logic [2:0] weight_6_30_reg;
logic [3:0] weight_6_31_reg;
logic [3:0] weight_6_32_reg;
logic [3:0] weight_6_33_reg;
logic [3:0] weight_6_34_reg;
logic [3:0] weight_6_35_reg;
logic [3:0] weight_6_36_reg;
logic [3:0] weight_6_37_reg;
logic [3:0] weight_6_38_reg;
logic [3:0] weight_6_39_reg;
logic [3:0] weight_6_40_reg;
logic [3:0] weight_6_41_reg;
logic [3:0] weight_6_42_reg;
logic [3:0] weight_6_43_reg;
logic [3:0] weight_6_44_reg;
logic [3:0] weight_6_45_reg;
logic [3:0] weight_6_46_reg;
logic [3:0] weight_6_47_reg;
logic [3:0] weight_6_48_reg;
logic [3:0] weight_6_49_reg;
logic [3:0] weight_6_50_reg;
logic [3:0] weight_6_51_reg;
logic [3:0] weight_6_52_reg;
logic [2:0] weight_6_53_reg;
logic [2:0] weight_6_54_reg;
logic [2:0] weight_6_55_reg;
logic [2:0] weight_6_56_reg;
logic [2:0] weight_6_57_reg;
logic [2:0] weight_6_58_reg;
logic [2:0] weight_6_59_reg;
logic [2:0] weight_6_60_reg;
logic [1:0] weight_6_61_reg;
logic [1:0] weight_6_62_reg;

// Second pipeline stage
always_ff @(posedge clk, negedge nrst) begin
    if (~nrst | multiplier_if.ready) begin
        en_reg_3 <= '0;
        weight_6_0_reg <= '0;
        weight_6_1_reg <= '0;
        weight_6_2_reg <= '0;
        weight_6_3_reg <= '0;
        weight_6_4_reg <= '0;
        weight_6_5_reg <= '0;
        weight_6_6_reg <= '0;
        weight_6_7_reg <= '0;
        weight_6_8_reg <= '0;
        weight_6_9_reg <= '0;
        weight_6_10_reg <= '0;
        weight_6_11_reg <= '0;
        weight_6_12_reg <= '0;
        weight_6_13_reg <= '0;
        weight_6_14_reg <= '0;
        weight_6_15_reg <= '0;
        weight_6_16_reg <= '0;
        weight_6_17_reg <= '0;
        weight_6_18_reg <= '0;
        weight_6_19_reg <= '0;
        weight_6_20_reg <= '0;
        weight_6_21_reg <= '0;
        weight_6_22_reg <= '0;
        weight_6_23_reg <= '0;
        weight_6_24_reg <= '0;
        weight_6_25_reg <= '0;
        weight_6_26_reg <= '0;
        weight_6_27_reg <= '0;
        weight_6_28_reg <= '0;
        weight_6_29_reg <= '0;
        weight_6_30_reg <= '0;
        weight_6_31_reg <= '0;
        weight_6_32_reg <= '0;
        weight_6_33_reg <= '0;
        weight_6_34_reg <= '0;
        weight_6_35_reg <= '0;
        weight_6_36_reg <= '0;
        weight_6_37_reg <= '0;
        weight_6_38_reg <= '0;
        weight_6_39_reg <= '0;
        weight_6_40_reg <= '0;
        weight_6_41_reg <= '0;
        weight_6_42_reg <= '0;
        weight_6_43_reg <= '0;
        weight_6_44_reg <= '0;
        weight_6_45_reg <= '0;
        weight_6_46_reg <= '0;
        weight_6_47_reg <= '0;
        weight_6_48_reg <= '0;
        weight_6_49_reg <= '0;
        weight_6_50_reg <= '0;
        weight_6_51_reg <= '0;
        weight_6_52_reg <= '0;
        weight_6_53_reg <= '0;
        weight_6_54_reg <= '0;
        weight_6_55_reg <= '0;
        weight_6_56_reg <= '0;
        weight_6_57_reg <= '0;
        weight_6_58_reg <= '0;
        weight_6_59_reg <= '0;
        weight_6_60_reg <= '0;
        weight_6_61_reg <= '0;
        weight_6_62_reg <= '0;
    end else begin
        en_reg_3 <= en_reg_2;
        weight_6_0_reg <= weight_6_0;
        weight_6_1_reg <= weight_6_1;
        weight_6_2_reg <= weight_6_2;
        weight_6_3_reg <= weight_6_3;
        weight_6_4_reg <= weight_6_4;
        weight_6_5_reg <= weight_6_5;
        weight_6_6_reg <= weight_6_6;
        weight_6_7_reg <= weight_6_7;
        weight_6_8_reg <= weight_6_8;
        weight_6_9_reg <= weight_6_9;
        weight_6_10_reg <= weight_6_10;
        weight_6_11_reg <= weight_6_11;
        weight_6_12_reg <= weight_6_12;
        weight_6_13_reg <= weight_6_13;
        weight_6_14_reg <= weight_6_14;
        weight_6_15_reg <= weight_6_15;
        weight_6_16_reg <= weight_6_16;
        weight_6_17_reg <= weight_6_17;
        weight_6_18_reg <= weight_6_18;
        weight_6_19_reg <= weight_6_19;
        weight_6_20_reg <= weight_6_20;
        weight_6_21_reg <= weight_6_21;
        weight_6_22_reg <= weight_6_22;
        weight_6_23_reg <= weight_6_23;
        weight_6_24_reg <= weight_6_24;
        weight_6_25_reg <= weight_6_25;
        weight_6_26_reg <= weight_6_26;
        weight_6_27_reg <= weight_6_27;
        weight_6_28_reg <= weight_6_28;
        weight_6_29_reg <= weight_6_29;
        weight_6_30_reg <= weight_6_30;
        weight_6_31_reg <= weight_6_31;
        weight_6_32_reg <= weight_6_32;
        weight_6_33_reg <= weight_6_33;
        weight_6_34_reg <= weight_6_34;
        weight_6_35_reg <= weight_6_35;
        weight_6_36_reg <= weight_6_36;
        weight_6_37_reg <= weight_6_37;
        weight_6_38_reg <= weight_6_38;
        weight_6_39_reg <= weight_6_39;
        weight_6_40_reg <= weight_6_40;
        weight_6_41_reg <= weight_6_41;
        weight_6_42_reg <= weight_6_42;
        weight_6_43_reg <= weight_6_43;
        weight_6_44_reg <= weight_6_44;
        weight_6_45_reg <= weight_6_45;
        weight_6_46_reg <= weight_6_46;
        weight_6_47_reg <= weight_6_47;
        weight_6_48_reg <= weight_6_48;
        weight_6_49_reg <= weight_6_49;
        weight_6_50_reg <= weight_6_50;
        weight_6_51_reg <= weight_6_51;
        weight_6_52_reg <= weight_6_52;
        weight_6_53_reg <= weight_6_53;
        weight_6_54_reg <= weight_6_54;
        weight_6_55_reg <= weight_6_55;
        weight_6_56_reg <= weight_6_56;
        weight_6_57_reg <= weight_6_57;
        weight_6_58_reg <= weight_6_58;
        weight_6_59_reg <= weight_6_59;
        weight_6_60_reg <= weight_6_60;
        weight_6_61_reg <= weight_6_61;
        weight_6_62_reg <= weight_6_62;
    end
end

assign weight_6_0 = weight_5_0;
assign weight_6_1 = weight_5_1;
assign weight_6_2 = weight_5_2;
assign weight_6_3 = weight_5_3;
assign weight_6_4 = weight_5_4;
assign weight_6_5 = weight_5_5;
half_adder ha94(.a(weight_5_6[0]), .b(weight_5_6[1]), .sum(weight_6_6), .cout(weight_6_7[0]));
half_adder ha95(.a(weight_5_7[0]), .b(weight_5_7[1]), .sum(weight_6_7[1]), .cout(weight_6_8[0]));
half_adder ha96(.a(weight_5_8[0]), .b(weight_5_8[1]), .sum(weight_6_8[1]), .cout(weight_6_9[0]));
half_adder ha97(.a(weight_5_9[0]), .b(weight_5_9[1]), .sum(weight_6_9[1]), .cout(weight_6_10[0]));
half_adder ha98(.a(weight_5_10[0]), .b(weight_5_10[1]), .sum(weight_6_10[1]), .cout(weight_6_11[0]));
half_adder ha99(.a(weight_5_11[0]), .b(weight_5_11[1]), .sum(weight_6_11[1]), .cout(weight_6_12[0]));
half_adder ha100(.a(weight_5_12[0]), .b(weight_5_12[1]), .sum(weight_6_12[1]), .cout(weight_6_13[0]));
half_adder ha101(.a(weight_5_13[0]), .b(weight_5_13[1]), .sum(weight_6_13[1]), .cout(weight_6_14[0]));
half_adder ha102(.a(weight_5_14[0]), .b(weight_5_14[1]), .sum(weight_6_14[1]), .cout(weight_6_15[0]));
full_adder fa813(.a(weight_5_15[0]), .b(weight_5_15[1]), .cin(weight_5_15[2]), .sum(weight_6_15[1]), .cout(weight_6_16[0]));
full_adder fa814(.a(weight_5_16[0]), .b(weight_5_16[1]), .cin(weight_5_16[2]), .sum(weight_6_16[1]), .cout(weight_6_17[0]));
full_adder fa815(.a(weight_5_17[0]), .b(weight_5_17[1]), .cin(weight_5_17[2]), .sum(weight_6_17[1]), .cout(weight_6_18[0]));
full_adder fa816(.a(weight_5_18[0]), .b(weight_5_18[1]), .cin(weight_5_18[2]), .sum(weight_6_18[1]), .cout(weight_6_19[0]));
full_adder fa817(.a(weight_5_19[0]), .b(weight_5_19[1]), .cin(weight_5_19[2]), .sum(weight_6_19[1]), .cout(weight_6_20[0]));
full_adder fa818(.a(weight_5_20[0]), .b(weight_5_20[1]), .cin(weight_5_20[2]), .sum(weight_6_20[1]), .cout(weight_6_21[0]));
full_adder fa819(.a(weight_5_21[0]), .b(weight_5_21[1]), .cin(weight_5_21[2]), .sum(weight_6_21[1]), .cout(weight_6_22[0]));
full_adder fa820(.a(weight_5_22[0]), .b(weight_5_22[1]), .cin(weight_5_22[2]), .sum(weight_6_22[1]), .cout(weight_6_23[0]));
full_adder fa821(.a(weight_5_23[0]), .b(weight_5_23[1]), .cin(weight_5_23[2]), .sum(weight_6_23[1]), .cout(weight_6_24[0]));
full_adder fa822(.a(weight_5_24[0]), .b(weight_5_24[1]), .cin(weight_5_24[2]), .sum(weight_6_24[1]), .cout(weight_6_25[0]));
full_adder fa823(.a(weight_5_25[0]), .b(weight_5_25[1]), .cin(weight_5_25[2]), .sum(weight_6_25[1]), .cout(weight_6_26[0]));
full_adder fa824(.a(weight_5_26[0]), .b(weight_5_26[1]), .cin(weight_5_26[2]), .sum(weight_6_26[1]), .cout(weight_6_27[0]));
full_adder fa825(.a(weight_5_27[0]), .b(weight_5_27[1]), .cin(weight_5_27[2]), .sum(weight_6_27[1]), .cout(weight_6_28[0]));
full_adder fa826(.a(weight_5_28[0]), .b(weight_5_28[1]), .cin(weight_5_28[2]), .sum(weight_6_28[1]), .cout(weight_6_29[0]));
full_adder fa827(.a(weight_5_29[0]), .b(weight_5_29[1]), .cin(weight_5_29[2]), .sum(weight_6_29[1]), .cout(weight_6_30[0]));
full_adder fa828(.a(weight_5_30[0]), .b(weight_5_30[1]), .cin(weight_5_30[2]), .sum(weight_6_30[1]), .cout(weight_6_31[0]));
full_adder fa829(.a(weight_5_31[0]), .b(weight_5_31[1]), .cin(weight_5_31[2]), .sum(weight_6_31[1]), .cout(weight_6_32[0]));
full_adder fa830(.a(weight_5_32[0]), .b(weight_5_32[1]), .cin(weight_5_32[2]), .sum(weight_6_32[1]), .cout(weight_6_33[0]));
full_adder fa831(.a(weight_5_33[0]), .b(weight_5_33[1]), .cin(weight_5_33[2]), .sum(weight_6_33[1]), .cout(weight_6_34[0]));
full_adder fa832(.a(weight_5_34[0]), .b(weight_5_34[1]), .cin(weight_5_34[2]), .sum(weight_6_34[1]), .cout(weight_6_35[0]));
full_adder fa833(.a(weight_5_35[0]), .b(weight_5_35[1]), .cin(weight_5_35[2]), .sum(weight_6_35[1]), .cout(weight_6_36[0]));
full_adder fa834(.a(weight_5_36[0]), .b(weight_5_36[1]), .cin(weight_5_36[2]), .sum(weight_6_36[1]), .cout(weight_6_37[0]));
full_adder fa835(.a(weight_5_37[0]), .b(weight_5_37[1]), .cin(weight_5_37[2]), .sum(weight_6_37[1]), .cout(weight_6_38[0]));
full_adder fa836(.a(weight_5_38[0]), .b(weight_5_38[1]), .cin(weight_5_38[2]), .sum(weight_6_38[1]), .cout(weight_6_39[0]));
full_adder fa837(.a(weight_5_39[0]), .b(weight_5_39[1]), .cin(weight_5_39[2]), .sum(weight_6_39[1]), .cout(weight_6_40[0]));
full_adder fa838(.a(weight_5_40[0]), .b(weight_5_40[1]), .cin(weight_5_40[2]), .sum(weight_6_40[1]), .cout(weight_6_41[0]));
full_adder fa839(.a(weight_5_41[0]), .b(weight_5_41[1]), .cin(weight_5_41[2]), .sum(weight_6_41[1]), .cout(weight_6_42[0]));
full_adder fa840(.a(weight_5_42[0]), .b(weight_5_42[1]), .cin(weight_5_42[2]), .sum(weight_6_42[1]), .cout(weight_6_43[0]));
full_adder fa841(.a(weight_5_43[0]), .b(weight_5_43[1]), .cin(weight_5_43[2]), .sum(weight_6_43[1]), .cout(weight_6_44[0]));
full_adder fa842(.a(weight_5_44[0]), .b(weight_5_44[1]), .cin(weight_5_44[2]), .sum(weight_6_44[1]), .cout(weight_6_45[0]));
full_adder fa843(.a(weight_5_45[0]), .b(weight_5_45[1]), .cin(weight_5_45[2]), .sum(weight_6_45[1]), .cout(weight_6_46[0]));
half_adder ha103(.a(weight_5_46[0]), .b(weight_5_46[1]), .sum(weight_6_46[1]), .cout(weight_6_47[0]));
half_adder ha104(.a(weight_5_47[0]), .b(weight_5_47[1]), .sum(weight_6_47[1]), .cout(weight_6_48[0]));
half_adder ha105(.a(weight_5_48[0]), .b(weight_5_48[1]), .sum(weight_6_48[1]), .cout(weight_6_49[0]));
half_adder ha106(.a(weight_5_49[0]), .b(weight_5_49[1]), .sum(weight_6_49[1]), .cout(weight_6_50[0]));
half_adder ha107(.a(weight_5_50[0]), .b(weight_5_50[1]), .sum(weight_6_50[1]), .cout(weight_6_51[0]));
half_adder ha108(.a(weight_5_51[0]), .b(weight_5_51[1]), .sum(weight_6_51[1]), .cout(weight_6_52[0]));
assign weight_6_52[1] = weight_5_52[0];
assign weight_6_53[0] = weight_5_53[0];
assign weight_6_54[0] = weight_5_54[0];
assign weight_6_55[0] = weight_5_55[0];
assign weight_6_56[0] = weight_5_56[0];
assign weight_6_57[0] = weight_5_57[0];
assign weight_6_58[0] = weight_5_58[0];
assign weight_6_59[0] = weight_5_59[0];
assign weight_6_60[0] = weight_5_60[0];
assign weight_6_22[2] = weight_5_22[3];
assign weight_6_23[2] = weight_5_23[3];
assign weight_6_24[2] = weight_5_24[3];
assign weight_6_25[2] = weight_5_25[3];
assign weight_6_26[2] = weight_5_26[3];
assign weight_6_27[2] = weight_5_27[3];
assign weight_6_28[2] = weight_5_28[3];
assign weight_6_29[2] = weight_5_29[3];
assign weight_6_30[2] = weight_5_30[3];
assign weight_6_31[2] = weight_5_31[3];
assign weight_6_32[2] = weight_5_32[3];
assign weight_6_33[2] = weight_5_33[3];
assign weight_6_34[2] = weight_5_34[3];
assign weight_6_35[2] = weight_5_35[3];
assign weight_6_36[2] = weight_5_36[3];
assign weight_6_37[2] = weight_5_37[3];
assign weight_6_38[2] = weight_5_38[3];
assign weight_6_39[2] = weight_5_39[3];
assign weight_6_40[2] = weight_5_40[3];
assign weight_6_41[2] = weight_5_41[3];
assign weight_6_42[2] = weight_5_42[3];
assign weight_6_43[2] = weight_5_43[3];
assign weight_6_44[2] = weight_5_44[3];
assign weight_6_45[2] = weight_5_45[3];
assign weight_6_46[2] = weight_5_46[2];
assign weight_6_47[2] = weight_5_47[2];
assign weight_6_48[2] = weight_5_48[2];
assign weight_6_49[2] = weight_5_49[2];
assign weight_6_50[2] = weight_5_50[2];
assign weight_6_51[2] = weight_5_51[2];
assign weight_6_52[2] = weight_5_52[1];
assign weight_6_53[1] = weight_5_53[1];
assign weight_6_54[1] = weight_5_54[1];
assign weight_6_55[1] = weight_5_55[1];
assign weight_6_56[1] = weight_5_56[1];
assign weight_6_57[1] = weight_5_57[1];
assign weight_6_58[1] = weight_5_58[1];
assign weight_6_59[1] = weight_5_59[1];
assign weight_6_60[1] = weight_5_60[1];
assign weight_6_61[0] = weight_5_61[0];
assign weight_6_62[0] = weight_5_62[0];
assign weight_6_31[3] = weight_5_31[4];
assign weight_6_32[3] = weight_5_32[4];
assign weight_6_33[3] = weight_5_33[4];
assign weight_6_34[3] = weight_5_34[4];
assign weight_6_35[3] = weight_5_35[4];
assign weight_6_36[3] = weight_5_36[4];
assign weight_6_37[3] = weight_5_37[4];
assign weight_6_38[3] = weight_5_38[4];
assign weight_6_39[3] = weight_5_39[4];
assign weight_6_40[3] = weight_5_40[4];
assign weight_6_41[3] = weight_5_41[4];
assign weight_6_42[3] = weight_5_42[4];
assign weight_6_43[3] = weight_5_43[4];
assign weight_6_44[3] = weight_5_44[4];
assign weight_6_45[3] = weight_5_45[4];
assign weight_6_46[3] = weight_5_46[3];
assign weight_6_47[3] = weight_5_47[3];
assign weight_6_48[3] = weight_5_48[3];
assign weight_6_49[3] = weight_5_49[3];
assign weight_6_50[3] = weight_5_50[3];
assign weight_6_51[3] = weight_5_51[3];
assign weight_6_52[3] = weight_5_52[2];
assign weight_6_53[2] = weight_5_53[2];
assign weight_6_54[2] = weight_5_54[2];
assign weight_6_55[2] = weight_5_55[2];
assign weight_6_56[2] = weight_5_56[2];
assign weight_6_57[2] = weight_5_57[2];
assign weight_6_58[2] = weight_5_58[2];
assign weight_6_59[2] = weight_5_59[2];
assign weight_6_60[2] = weight_5_60[2];
assign weight_6_61[1] = weight_5_61[1];
assign weight_6_62[1] = weight_5_62[1];
logic weight_7_0;
logic weight_7_1;
logic weight_7_2;
logic weight_7_3;
logic weight_7_4;
logic weight_7_5;
logic weight_7_6;
logic weight_7_7;
logic [1:0] weight_7_8;
logic [1:0] weight_7_9;
logic [1:0] weight_7_10;
logic [1:0] weight_7_11;
logic [1:0] weight_7_12;
logic [1:0] weight_7_13;
logic [1:0] weight_7_14;
logic [1:0] weight_7_15;
logic [1:0] weight_7_16;
logic [1:0] weight_7_17;
logic [1:0] weight_7_18;
logic [1:0] weight_7_19;
logic [1:0] weight_7_20;
logic [1:0] weight_7_21;
logic [1:0] weight_7_22;
logic [1:0] weight_7_23;
logic [1:0] weight_7_24;
logic [1:0] weight_7_25;
logic [1:0] weight_7_26;
logic [1:0] weight_7_27;
logic [1:0] weight_7_28;
logic [1:0] weight_7_29;
logic [1:0] weight_7_30;
logic [2:0] weight_7_31;
logic [2:0] weight_7_32;
logic [2:0] weight_7_33;
logic [2:0] weight_7_34;
logic [2:0] weight_7_35;
logic [2:0] weight_7_36;
logic [2:0] weight_7_37;
logic [2:0] weight_7_38;
logic [2:0] weight_7_39;
logic [2:0] weight_7_40;
logic [2:0] weight_7_41;
logic [2:0] weight_7_42;
logic [2:0] weight_7_43;
logic [2:0] weight_7_44;
logic [2:0] weight_7_45;
logic [2:0] weight_7_46;
logic [2:0] weight_7_47;
logic [2:0] weight_7_48;
logic [2:0] weight_7_49;
logic [2:0] weight_7_50;
logic [2:0] weight_7_51;
logic [2:0] weight_7_52;
logic [2:0] weight_7_53;
logic [2:0] weight_7_54;
logic [2:0] weight_7_55;
logic [2:0] weight_7_56;
logic [2:0] weight_7_57;
logic [2:0] weight_7_58;
logic [2:0] weight_7_59;
logic [2:0] weight_7_60;
logic [2:0] weight_7_61;
logic [1:0] weight_7_62;
assign weight_7_0 = weight_6_0_reg;
assign weight_7_1 = weight_6_1_reg;
assign weight_7_2 = weight_6_2_reg;
assign weight_7_3 = weight_6_3_reg;
assign weight_7_4 = weight_6_4_reg;
assign weight_7_5 = weight_6_5_reg;
assign weight_7_6 = weight_6_6_reg;
half_adder ha109(.a(weight_6_7_reg[0]), .b(weight_6_7_reg[1]), .sum(weight_7_7), .cout(weight_7_8[0]));
half_adder ha110(.a(weight_6_8_reg[0]), .b(weight_6_8_reg[1]), .sum(weight_7_8[1]), .cout(weight_7_9[0]));
half_adder ha111(.a(weight_6_9_reg[0]), .b(weight_6_9_reg[1]), .sum(weight_7_9[1]), .cout(weight_7_10[0]));
half_adder ha112(.a(weight_6_10_reg[0]), .b(weight_6_10_reg[1]), .sum(weight_7_10[1]), .cout(weight_7_11[0]));
half_adder ha113(.a(weight_6_11_reg[0]), .b(weight_6_11_reg[1]), .sum(weight_7_11[1]), .cout(weight_7_12[0]));
half_adder ha114(.a(weight_6_12_reg[0]), .b(weight_6_12_reg[1]), .sum(weight_7_12[1]), .cout(weight_7_13[0]));
half_adder ha115(.a(weight_6_13_reg[0]), .b(weight_6_13_reg[1]), .sum(weight_7_13[1]), .cout(weight_7_14[0]));
half_adder ha116(.a(weight_6_14_reg[0]), .b(weight_6_14_reg[1]), .sum(weight_7_14[1]), .cout(weight_7_15[0]));
half_adder ha117(.a(weight_6_15_reg[0]), .b(weight_6_15_reg[1]), .sum(weight_7_15[1]), .cout(weight_7_16[0]));
half_adder ha118(.a(weight_6_16_reg[0]), .b(weight_6_16_reg[1]), .sum(weight_7_16[1]), .cout(weight_7_17[0]));
half_adder ha119(.a(weight_6_17_reg[0]), .b(weight_6_17_reg[1]), .sum(weight_7_17[1]), .cout(weight_7_18[0]));
half_adder ha120(.a(weight_6_18_reg[0]), .b(weight_6_18_reg[1]), .sum(weight_7_18[1]), .cout(weight_7_19[0]));
half_adder ha121(.a(weight_6_19_reg[0]), .b(weight_6_19_reg[1]), .sum(weight_7_19[1]), .cout(weight_7_20[0]));
half_adder ha122(.a(weight_6_20_reg[0]), .b(weight_6_20_reg[1]), .sum(weight_7_20[1]), .cout(weight_7_21[0]));
half_adder ha123(.a(weight_6_21_reg[0]), .b(weight_6_21_reg[1]), .sum(weight_7_21[1]), .cout(weight_7_22[0]));
full_adder fa844(.a(weight_6_22_reg[0]), .b(weight_6_22_reg[1]), .cin(weight_6_22_reg[2]), .sum(weight_7_22[1]), .cout(weight_7_23[0]));
full_adder fa845(.a(weight_6_23_reg[0]), .b(weight_6_23_reg[1]), .cin(weight_6_23_reg[2]), .sum(weight_7_23[1]), .cout(weight_7_24[0]));
full_adder fa846(.a(weight_6_24_reg[0]), .b(weight_6_24_reg[1]), .cin(weight_6_24_reg[2]), .sum(weight_7_24[1]), .cout(weight_7_25[0]));
full_adder fa847(.a(weight_6_25_reg[0]), .b(weight_6_25_reg[1]), .cin(weight_6_25_reg[2]), .sum(weight_7_25[1]), .cout(weight_7_26[0]));
full_adder fa848(.a(weight_6_26_reg[0]), .b(weight_6_26_reg[1]), .cin(weight_6_26_reg[2]), .sum(weight_7_26[1]), .cout(weight_7_27[0]));
full_adder fa849(.a(weight_6_27_reg[0]), .b(weight_6_27_reg[1]), .cin(weight_6_27_reg[2]), .sum(weight_7_27[1]), .cout(weight_7_28[0]));
full_adder fa850(.a(weight_6_28_reg[0]), .b(weight_6_28_reg[1]), .cin(weight_6_28_reg[2]), .sum(weight_7_28[1]), .cout(weight_7_29[0]));
full_adder fa851(.a(weight_6_29_reg[0]), .b(weight_6_29_reg[1]), .cin(weight_6_29_reg[2]), .sum(weight_7_29[1]), .cout(weight_7_30[0]));
full_adder fa852(.a(weight_6_30_reg[0]), .b(weight_6_30_reg[1]), .cin(weight_6_30_reg[2]), .sum(weight_7_30[1]), .cout(weight_7_31[0]));
full_adder fa853(.a(weight_6_31_reg[0]), .b(weight_6_31_reg[1]), .cin(weight_6_31_reg[2]), .sum(weight_7_31[1]), .cout(weight_7_32[0]));
full_adder fa854(.a(weight_6_32_reg[0]), .b(weight_6_32_reg[1]), .cin(weight_6_32_reg[2]), .sum(weight_7_32[1]), .cout(weight_7_33[0]));
full_adder fa855(.a(weight_6_33_reg[0]), .b(weight_6_33_reg[1]), .cin(weight_6_33_reg[2]), .sum(weight_7_33[1]), .cout(weight_7_34[0]));
full_adder fa856(.a(weight_6_34_reg[0]), .b(weight_6_34_reg[1]), .cin(weight_6_34_reg[2]), .sum(weight_7_34[1]), .cout(weight_7_35[0]));
full_adder fa857(.a(weight_6_35_reg[0]), .b(weight_6_35_reg[1]), .cin(weight_6_35_reg[2]), .sum(weight_7_35[1]), .cout(weight_7_36[0]));
full_adder fa858(.a(weight_6_36_reg[0]), .b(weight_6_36_reg[1]), .cin(weight_6_36_reg[2]), .sum(weight_7_36[1]), .cout(weight_7_37[0]));
full_adder fa859(.a(weight_6_37_reg[0]), .b(weight_6_37_reg[1]), .cin(weight_6_37_reg[2]), .sum(weight_7_37[1]), .cout(weight_7_38[0]));
full_adder fa860(.a(weight_6_38_reg[0]), .b(weight_6_38_reg[1]), .cin(weight_6_38_reg[2]), .sum(weight_7_38[1]), .cout(weight_7_39[0]));
full_adder fa861(.a(weight_6_39_reg[0]), .b(weight_6_39_reg[1]), .cin(weight_6_39_reg[2]), .sum(weight_7_39[1]), .cout(weight_7_40[0]));
full_adder fa862(.a(weight_6_40_reg[0]), .b(weight_6_40_reg[1]), .cin(weight_6_40_reg[2]), .sum(weight_7_40[1]), .cout(weight_7_41[0]));
full_adder fa863(.a(weight_6_41_reg[0]), .b(weight_6_41_reg[1]), .cin(weight_6_41_reg[2]), .sum(weight_7_41[1]), .cout(weight_7_42[0]));
full_adder fa864(.a(weight_6_42_reg[0]), .b(weight_6_42_reg[1]), .cin(weight_6_42_reg[2]), .sum(weight_7_42[1]), .cout(weight_7_43[0]));
full_adder fa865(.a(weight_6_43_reg[0]), .b(weight_6_43_reg[1]), .cin(weight_6_43_reg[2]), .sum(weight_7_43[1]), .cout(weight_7_44[0]));
full_adder fa866(.a(weight_6_44_reg[0]), .b(weight_6_44_reg[1]), .cin(weight_6_44_reg[2]), .sum(weight_7_44[1]), .cout(weight_7_45[0]));
full_adder fa867(.a(weight_6_45_reg[0]), .b(weight_6_45_reg[1]), .cin(weight_6_45_reg[2]), .sum(weight_7_45[1]), .cout(weight_7_46[0]));
full_adder fa868(.a(weight_6_46_reg[0]), .b(weight_6_46_reg[1]), .cin(weight_6_46_reg[2]), .sum(weight_7_46[1]), .cout(weight_7_47[0]));
full_adder fa869(.a(weight_6_47_reg[0]), .b(weight_6_47_reg[1]), .cin(weight_6_47_reg[2]), .sum(weight_7_47[1]), .cout(weight_7_48[0]));
full_adder fa870(.a(weight_6_48_reg[0]), .b(weight_6_48_reg[1]), .cin(weight_6_48_reg[2]), .sum(weight_7_48[1]), .cout(weight_7_49[0]));
full_adder fa871(.a(weight_6_49_reg[0]), .b(weight_6_49_reg[1]), .cin(weight_6_49_reg[2]), .sum(weight_7_49[1]), .cout(weight_7_50[0]));
full_adder fa872(.a(weight_6_50_reg[0]), .b(weight_6_50_reg[1]), .cin(weight_6_50_reg[2]), .sum(weight_7_50[1]), .cout(weight_7_51[0]));
full_adder fa873(.a(weight_6_51_reg[0]), .b(weight_6_51_reg[1]), .cin(weight_6_51_reg[2]), .sum(weight_7_51[1]), .cout(weight_7_52[0]));
full_adder fa874(.a(weight_6_52_reg[0]), .b(weight_6_52_reg[1]), .cin(weight_6_52_reg[2]), .sum(weight_7_52[1]), .cout(weight_7_53[0]));
half_adder ha124(.a(weight_6_53_reg[0]), .b(weight_6_53_reg[1]), .sum(weight_7_53[1]), .cout(weight_7_54[0]));
half_adder ha125(.a(weight_6_54_reg[0]), .b(weight_6_54_reg[1]), .sum(weight_7_54[1]), .cout(weight_7_55[0]));
half_adder ha126(.a(weight_6_55_reg[0]), .b(weight_6_55_reg[1]), .sum(weight_7_55[1]), .cout(weight_7_56[0]));
half_adder ha127(.a(weight_6_56_reg[0]), .b(weight_6_56_reg[1]), .sum(weight_7_56[1]), .cout(weight_7_57[0]));
half_adder ha128(.a(weight_6_57_reg[0]), .b(weight_6_57_reg[1]), .sum(weight_7_57[1]), .cout(weight_7_58[0]));
half_adder ha129(.a(weight_6_58_reg[0]), .b(weight_6_58_reg[1]), .sum(weight_7_58[1]), .cout(weight_7_59[0]));
half_adder ha130(.a(weight_6_59_reg[0]), .b(weight_6_59_reg[1]), .sum(weight_7_59[1]), .cout(weight_7_60[0]));
half_adder ha131(.a(weight_6_60_reg[0]), .b(weight_6_60_reg[1]), .sum(weight_7_60[1]), .cout(weight_7_61[0]));
assign weight_7_61[1] = weight_6_61_reg[0];
assign weight_7_62[0] = weight_6_62_reg[0];
assign weight_7_31[2] = weight_6_31_reg[3];
assign weight_7_32[2] = weight_6_32_reg[3];
assign weight_7_33[2] = weight_6_33_reg[3];
assign weight_7_34[2] = weight_6_34_reg[3];
assign weight_7_35[2] = weight_6_35_reg[3];
assign weight_7_36[2] = weight_6_36_reg[3];
assign weight_7_37[2] = weight_6_37_reg[3];
assign weight_7_38[2] = weight_6_38_reg[3];
assign weight_7_39[2] = weight_6_39_reg[3];
assign weight_7_40[2] = weight_6_40_reg[3];
assign weight_7_41[2] = weight_6_41_reg[3];
assign weight_7_42[2] = weight_6_42_reg[3];
assign weight_7_43[2] = weight_6_43_reg[3];
assign weight_7_44[2] = weight_6_44_reg[3];
assign weight_7_45[2] = weight_6_45_reg[3];
assign weight_7_46[2] = weight_6_46_reg[3];
assign weight_7_47[2] = weight_6_47_reg[3];
assign weight_7_48[2] = weight_6_48_reg[3];
assign weight_7_49[2] = weight_6_49_reg[3];
assign weight_7_50[2] = weight_6_50_reg[3];
assign weight_7_51[2] = weight_6_51_reg[3];
assign weight_7_52[2] = weight_6_52_reg[3];
assign weight_7_53[2] = weight_6_53_reg[2];
assign weight_7_54[2] = weight_6_54_reg[2];
assign weight_7_55[2] = weight_6_55_reg[2];
assign weight_7_56[2] = weight_6_56_reg[2];
assign weight_7_57[2] = weight_6_57_reg[2];
assign weight_7_58[2] = weight_6_58_reg[2];
assign weight_7_59[2] = weight_6_59_reg[2];
assign weight_7_60[2] = weight_6_60_reg[2];
assign weight_7_61[2] = weight_6_61_reg[1];
assign weight_7_62[1] = weight_6_62_reg[1];
logic weight_8_0;
logic weight_8_1;
logic weight_8_2;
logic weight_8_3;
logic weight_8_4;
logic weight_8_5;
logic weight_8_6;
logic weight_8_7;
logic weight_8_8;
logic [1:0] weight_8_9;
logic [1:0] weight_8_10;
logic [1:0] weight_8_11;
logic [1:0] weight_8_12;
logic [1:0] weight_8_13;
logic [1:0] weight_8_14;
logic [1:0] weight_8_15;
logic [1:0] weight_8_16;
logic [1:0] weight_8_17;
logic [1:0] weight_8_18;
logic [1:0] weight_8_19;
logic [1:0] weight_8_20;
logic [1:0] weight_8_21;
logic [1:0] weight_8_22;
logic [1:0] weight_8_23;
logic [1:0] weight_8_24;
logic [1:0] weight_8_25;
logic [1:0] weight_8_26;
logic [1:0] weight_8_27;
logic [1:0] weight_8_28;
logic [1:0] weight_8_29;
logic [1:0] weight_8_30;
logic [1:0] weight_8_31;
logic [1:0] weight_8_32;
logic [1:0] weight_8_33;
logic [1:0] weight_8_34;
logic [1:0] weight_8_35;
logic [1:0] weight_8_36;
logic [1:0] weight_8_37;
logic [1:0] weight_8_38;
logic [1:0] weight_8_39;
logic [1:0] weight_8_40;
logic [1:0] weight_8_41;
logic [1:0] weight_8_42;
logic [1:0] weight_8_43;
logic [1:0] weight_8_44;
logic [1:0] weight_8_45;
logic [1:0] weight_8_46;
logic [1:0] weight_8_47;
logic [1:0] weight_8_48;
logic [1:0] weight_8_49;
logic [1:0] weight_8_50;
logic [1:0] weight_8_51;
logic [1:0] weight_8_52;
logic [1:0] weight_8_53;
logic [1:0] weight_8_54;
logic [1:0] weight_8_55;
logic [1:0] weight_8_56;
logic [1:0] weight_8_57;
logic [1:0] weight_8_58;
logic [1:0] weight_8_59;
logic [1:0] weight_8_60;
logic [1:0] weight_8_61;
logic [1:0] weight_8_62;
logic weight_8_63;
assign weight_8_0 = weight_7_0;
assign weight_8_1 = weight_7_1;
assign weight_8_2 = weight_7_2;
assign weight_8_3 = weight_7_3;
assign weight_8_4 = weight_7_4;
assign weight_8_5 = weight_7_5;
assign weight_8_6 = weight_7_6;
assign weight_8_7 = weight_7_7;
half_adder ha132(.a(weight_7_8[0]), .b(weight_7_8[1]), .sum(weight_8_8), .cout(weight_8_9[0]));
half_adder ha133(.a(weight_7_9[0]), .b(weight_7_9[1]), .sum(weight_8_9[1]), .cout(weight_8_10[0]));
half_adder ha134(.a(weight_7_10[0]), .b(weight_7_10[1]), .sum(weight_8_10[1]), .cout(weight_8_11[0]));
half_adder ha135(.a(weight_7_11[0]), .b(weight_7_11[1]), .sum(weight_8_11[1]), .cout(weight_8_12[0]));
half_adder ha136(.a(weight_7_12[0]), .b(weight_7_12[1]), .sum(weight_8_12[1]), .cout(weight_8_13[0]));
half_adder ha137(.a(weight_7_13[0]), .b(weight_7_13[1]), .sum(weight_8_13[1]), .cout(weight_8_14[0]));
half_adder ha138(.a(weight_7_14[0]), .b(weight_7_14[1]), .sum(weight_8_14[1]), .cout(weight_8_15[0]));
half_adder ha139(.a(weight_7_15[0]), .b(weight_7_15[1]), .sum(weight_8_15[1]), .cout(weight_8_16[0]));
half_adder ha140(.a(weight_7_16[0]), .b(weight_7_16[1]), .sum(weight_8_16[1]), .cout(weight_8_17[0]));
half_adder ha141(.a(weight_7_17[0]), .b(weight_7_17[1]), .sum(weight_8_17[1]), .cout(weight_8_18[0]));
half_adder ha142(.a(weight_7_18[0]), .b(weight_7_18[1]), .sum(weight_8_18[1]), .cout(weight_8_19[0]));
half_adder ha143(.a(weight_7_19[0]), .b(weight_7_19[1]), .sum(weight_8_19[1]), .cout(weight_8_20[0]));
half_adder ha144(.a(weight_7_20[0]), .b(weight_7_20[1]), .sum(weight_8_20[1]), .cout(weight_8_21[0]));
half_adder ha145(.a(weight_7_21[0]), .b(weight_7_21[1]), .sum(weight_8_21[1]), .cout(weight_8_22[0]));
half_adder ha146(.a(weight_7_22[0]), .b(weight_7_22[1]), .sum(weight_8_22[1]), .cout(weight_8_23[0]));
half_adder ha147(.a(weight_7_23[0]), .b(weight_7_23[1]), .sum(weight_8_23[1]), .cout(weight_8_24[0]));
half_adder ha148(.a(weight_7_24[0]), .b(weight_7_24[1]), .sum(weight_8_24[1]), .cout(weight_8_25[0]));
half_adder ha149(.a(weight_7_25[0]), .b(weight_7_25[1]), .sum(weight_8_25[1]), .cout(weight_8_26[0]));
half_adder ha150(.a(weight_7_26[0]), .b(weight_7_26[1]), .sum(weight_8_26[1]), .cout(weight_8_27[0]));
half_adder ha151(.a(weight_7_27[0]), .b(weight_7_27[1]), .sum(weight_8_27[1]), .cout(weight_8_28[0]));
half_adder ha152(.a(weight_7_28[0]), .b(weight_7_28[1]), .sum(weight_8_28[1]), .cout(weight_8_29[0]));
half_adder ha153(.a(weight_7_29[0]), .b(weight_7_29[1]), .sum(weight_8_29[1]), .cout(weight_8_30[0]));
half_adder ha154(.a(weight_7_30[0]), .b(weight_7_30[1]), .sum(weight_8_30[1]), .cout(weight_8_31[0]));
full_adder fa875(.a(weight_7_31[0]), .b(weight_7_31[1]), .cin(weight_7_31[2]), .sum(weight_8_31[1]), .cout(weight_8_32[0]));
full_adder fa876(.a(weight_7_32[0]), .b(weight_7_32[1]), .cin(weight_7_32[2]), .sum(weight_8_32[1]), .cout(weight_8_33[0]));
full_adder fa877(.a(weight_7_33[0]), .b(weight_7_33[1]), .cin(weight_7_33[2]), .sum(weight_8_33[1]), .cout(weight_8_34[0]));
full_adder fa878(.a(weight_7_34[0]), .b(weight_7_34[1]), .cin(weight_7_34[2]), .sum(weight_8_34[1]), .cout(weight_8_35[0]));
full_adder fa879(.a(weight_7_35[0]), .b(weight_7_35[1]), .cin(weight_7_35[2]), .sum(weight_8_35[1]), .cout(weight_8_36[0]));
full_adder fa880(.a(weight_7_36[0]), .b(weight_7_36[1]), .cin(weight_7_36[2]), .sum(weight_8_36[1]), .cout(weight_8_37[0]));
full_adder fa881(.a(weight_7_37[0]), .b(weight_7_37[1]), .cin(weight_7_37[2]), .sum(weight_8_37[1]), .cout(weight_8_38[0]));
full_adder fa882(.a(weight_7_38[0]), .b(weight_7_38[1]), .cin(weight_7_38[2]), .sum(weight_8_38[1]), .cout(weight_8_39[0]));
full_adder fa883(.a(weight_7_39[0]), .b(weight_7_39[1]), .cin(weight_7_39[2]), .sum(weight_8_39[1]), .cout(weight_8_40[0]));
full_adder fa884(.a(weight_7_40[0]), .b(weight_7_40[1]), .cin(weight_7_40[2]), .sum(weight_8_40[1]), .cout(weight_8_41[0]));
full_adder fa885(.a(weight_7_41[0]), .b(weight_7_41[1]), .cin(weight_7_41[2]), .sum(weight_8_41[1]), .cout(weight_8_42[0]));
full_adder fa886(.a(weight_7_42[0]), .b(weight_7_42[1]), .cin(weight_7_42[2]), .sum(weight_8_42[1]), .cout(weight_8_43[0]));
full_adder fa887(.a(weight_7_43[0]), .b(weight_7_43[1]), .cin(weight_7_43[2]), .sum(weight_8_43[1]), .cout(weight_8_44[0]));
full_adder fa888(.a(weight_7_44[0]), .b(weight_7_44[1]), .cin(weight_7_44[2]), .sum(weight_8_44[1]), .cout(weight_8_45[0]));
full_adder fa889(.a(weight_7_45[0]), .b(weight_7_45[1]), .cin(weight_7_45[2]), .sum(weight_8_45[1]), .cout(weight_8_46[0]));
full_adder fa890(.a(weight_7_46[0]), .b(weight_7_46[1]), .cin(weight_7_46[2]), .sum(weight_8_46[1]), .cout(weight_8_47[0]));
full_adder fa891(.a(weight_7_47[0]), .b(weight_7_47[1]), .cin(weight_7_47[2]), .sum(weight_8_47[1]), .cout(weight_8_48[0]));
full_adder fa892(.a(weight_7_48[0]), .b(weight_7_48[1]), .cin(weight_7_48[2]), .sum(weight_8_48[1]), .cout(weight_8_49[0]));
full_adder fa893(.a(weight_7_49[0]), .b(weight_7_49[1]), .cin(weight_7_49[2]), .sum(weight_8_49[1]), .cout(weight_8_50[0]));
full_adder fa894(.a(weight_7_50[0]), .b(weight_7_50[1]), .cin(weight_7_50[2]), .sum(weight_8_50[1]), .cout(weight_8_51[0]));
full_adder fa895(.a(weight_7_51[0]), .b(weight_7_51[1]), .cin(weight_7_51[2]), .sum(weight_8_51[1]), .cout(weight_8_52[0]));
full_adder fa896(.a(weight_7_52[0]), .b(weight_7_52[1]), .cin(weight_7_52[2]), .sum(weight_8_52[1]), .cout(weight_8_53[0]));
full_adder fa897(.a(weight_7_53[0]), .b(weight_7_53[1]), .cin(weight_7_53[2]), .sum(weight_8_53[1]), .cout(weight_8_54[0]));
full_adder fa898(.a(weight_7_54[0]), .b(weight_7_54[1]), .cin(weight_7_54[2]), .sum(weight_8_54[1]), .cout(weight_8_55[0]));
full_adder fa899(.a(weight_7_55[0]), .b(weight_7_55[1]), .cin(weight_7_55[2]), .sum(weight_8_55[1]), .cout(weight_8_56[0]));
full_adder fa900(.a(weight_7_56[0]), .b(weight_7_56[1]), .cin(weight_7_56[2]), .sum(weight_8_56[1]), .cout(weight_8_57[0]));
full_adder fa901(.a(weight_7_57[0]), .b(weight_7_57[1]), .cin(weight_7_57[2]), .sum(weight_8_57[1]), .cout(weight_8_58[0]));
full_adder fa902(.a(weight_7_58[0]), .b(weight_7_58[1]), .cin(weight_7_58[2]), .sum(weight_8_58[1]), .cout(weight_8_59[0]));
full_adder fa903(.a(weight_7_59[0]), .b(weight_7_59[1]), .cin(weight_7_59[2]), .sum(weight_8_59[1]), .cout(weight_8_60[0]));
full_adder fa904(.a(weight_7_60[0]), .b(weight_7_60[1]), .cin(weight_7_60[2]), .sum(weight_8_60[1]), .cout(weight_8_61[0]));
full_adder fa905(.a(weight_7_61[0]), .b(weight_7_61[1]), .cin(weight_7_61[2]), .sum(weight_8_61[1]), .cout(weight_8_62[0]));
half_adder ha155(.a(weight_7_62[0]), .b(weight_7_62[1]), .sum(weight_8_62[1]), .cout(weight_8_63));
logic [63:0] final_sum_a;
logic [63:0] final_sum_b;
assign final_sum_a = {weight_8_63, weight_8_62[0], weight_8_61[0], weight_8_60[0], weight_8_59[0], weight_8_58[0], weight_8_57[0], weight_8_56[0], weight_8_55[0], weight_8_54[0], weight_8_53[0], weight_8_52[0], weight_8_51[0], weight_8_50[0], weight_8_49[0], weight_8_48[0], weight_8_47[0], weight_8_46[0], weight_8_45[0], weight_8_44[0], weight_8_43[0], weight_8_42[0], weight_8_41[0], weight_8_40[0], weight_8_39[0], weight_8_38[0], weight_8_37[0], weight_8_36[0], weight_8_35[0], weight_8_34[0], weight_8_33[0], weight_8_32[0], weight_8_31[0], weight_8_30[0], weight_8_29[0], weight_8_28[0], weight_8_27[0], weight_8_26[0], weight_8_25[0], weight_8_24[0], weight_8_23[0], weight_8_22[0], weight_8_21[0], weight_8_20[0], weight_8_19[0], weight_8_18[0], weight_8_17[0], weight_8_16[0], weight_8_15[0], weight_8_14[0], weight_8_13[0], weight_8_12[0], weight_8_11[0], weight_8_10[0], weight_8_9[0], weight_8_8, weight_8_7, weight_8_6, weight_8_5, weight_8_4, weight_8_3, weight_8_2, weight_8_1, weight_8_0};
assign final_sum_b = {1'b0, weight_8_62[1], weight_8_61[1], weight_8_60[1], weight_8_59[1], weight_8_58[1], weight_8_57[1], weight_8_56[1], weight_8_55[1], weight_8_54[1], weight_8_53[1], weight_8_52[1], weight_8_51[1], weight_8_50[1], weight_8_49[1], weight_8_48[1], weight_8_47[1], weight_8_46[1], weight_8_45[1], weight_8_44[1], weight_8_43[1], weight_8_42[1], weight_8_41[1], weight_8_40[1], weight_8_39[1], weight_8_38[1], weight_8_37[1], weight_8_36[1], weight_8_35[1], weight_8_34[1], weight_8_33[1], weight_8_32[1], weight_8_31[1], weight_8_30[1], weight_8_29[1], weight_8_28[1], weight_8_27[1], weight_8_26[1], weight_8_25[1], weight_8_24[1], weight_8_23[1], weight_8_22[1], weight_8_21[1], weight_8_20[1], weight_8_19[1], weight_8_18[1], weight_8_17[1], weight_8_16[1], weight_8_15[1], weight_8_14[1], weight_8_13[1], weight_8_12[1], weight_8_11[1], weight_8_10[1], weight_8_9[1], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};


always_comb begin
    multiplier_if.out = final_sum_a + final_sum_b;
    multiplier_if.ready = multiplier_if.en & en_reg_3;
    if(multiplier_if.is_signed_a && multiplier_if.is_signed_b) begin
        // If the signs are different, the result is negative
        if(multiplier_if.a[31] ^ multiplier_if.b[31]) begin
            multiplier_if.out = ~multiplier_if.out + 1;
        end
    end else if (multiplier_if.is_signed_a) begin
        // If the first number is negative, the result is negative
        if(multiplier_if.a[31]) begin
            multiplier_if.out = ~multiplier_if.out + 1;
        end
    end else if (multiplier_if.is_signed_b) begin
        // If the second number is negative, the result is negative
        if(multiplier_if.b[31]) begin
            multiplier_if.out = ~multiplier_if.out + 1;
        end
    end
end

endmodule